`timescale 1ns / 1ps

module pingpang
(
    input  wire        sys_clk ,      // ϵͳʱ�� 50MHz
    input  wire        sys_rst_n ,    // ��λ (����Ч)
    
    // ------------------------------------------
    // ���νӿ� (��������)
    // ------------------------------------------
    input  wire        data_en ,      // ���� Valid
    input  wire [63:0] data_in ,      // ���� Data
    output wire        o_upstream_ready, // ����������� Ready (��ѹ����)

    // ------------------------------------------
    // ���νӿ� (��������)
    // ------------------------------------------
    input  wire        i_downstream_ready, // ������������ Ready (���շ�ѹ)
    output wire        o_downstream_valid, // ����������� Valid
    output wire [63:0] data_out            // ��� Data
);

    //================================================
    // Internal Signals
    //================================================
    wire clk_50m ;
    wire rst_n ;

    // RAM1 �����ź�
    wire [63:0] ram1_rd_data ;
    wire [63:0] ram1_wr_data ;
    wire ram1_wr_en ;
    wire ram1_rd_en ;
    wire [5:0] ram1_wr_addr ;
    wire [5:0] ram1_rd_addr ;

    // RAM2 �����ź�
    wire [63:0] ram2_rd_data ;
    wire [63:0] ram2_wr_data ;
    wire ram2_wr_en ;
    wire ram2_rd_en ;
    wire [5:0] ram2_wr_addr ;
    wire [5:0] ram2_rd_addr ;

    // �򵥸�ֵ
    assign rst_n   = sys_rst_n ;
    assign clk_50m = sys_clk ;

    //================================================
    // 1. ʵ�������ƺ��� (ram_ctrl)
    //================================================
    ram_ctrl1 ram_ctrl_inst
    (
        .clk_50m      (clk_50m),
        .rst_n        (rst_n),
        
        // RAM ����ͨ·
        .ram1_rd_data (ram1_rd_data),
        .ram2_rd_data (ram2_rd_data),
        .ram1_wr_data (ram1_wr_data),
        .ram2_wr_data (ram2_wr_data),
        
        // RAM �����ź�
        .ram1_wr_en   (ram1_wr_en),
        .ram1_rd_en   (ram1_rd_en),
        .ram1_wr_addr (ram1_wr_addr),
        .ram1_rd_addr (ram1_rd_addr),
        
        .ram2_wr_en   (ram2_wr_en),
        .ram2_rd_en   (ram2_rd_en),
        .ram2_wr_addr (ram2_wr_addr),
        .ram2_rd_addr (ram2_rd_addr),

        // ��������
        .data_en          (data_en),
        .data_in          (data_in),
        .o_upstream_ready (o_upstream_ready), // ���������˿�
        
        // ��������
        .i_downstream_ready (i_downstream_ready), // ���������˿�
        .o_data_valid       (o_downstream_valid), // ���������˿�
        .data_out           (data_out)
    );

    //================================================
    // 2. ʵ���� RAM IP ��
    //================================================
    
    // RAM 1
    dist_mem_gen_0 sdp_ram1 (
        .clk (clk_50m),       // ����Ҫ������ʱ������
        .we  (ram1_wr_en),
        .a   (ram1_wr_addr),
        .d   (ram1_wr_data),
        .dpra(ram1_rd_addr),
        .dpo (ram1_rd_data)
    );

    // RAM 2
    dist_mem_gen_0 sdp_ram2 (
        .clk (clk_50m),       // ����Ҫ������ʱ������
        .we  (ram2_wr_en),
        .a   (ram2_wr_addr),
        .d   (ram2_wr_data),
        .dpra(ram2_rd_addr),
        .dpo (ram2_rd_data)
    );

endmodule