`timescale 1ns / 1ps
module ram_ctrl1
(
    input  wire        clk_50m ,
    input  wire        rst_n ,
    
    input  wire [63:0] ram1_rd_data, 
    input  wire [63:0] ram2_rd_data, 
    output wire [63:0] ram1_wr_data, 
    output wire [63:0] ram2_wr_data, 
    
    output reg         ram1_wr_en , 
    output reg         ram1_rd_en , 
    
    // 依然使用 7 位宽地址，确保能计数�? 64
    output reg  [6:0]  ram1_wr_addr, 
    output reg  [5:0]  ram1_rd_addr, 
    
    output reg         ram2_wr_en , 
    output reg         ram2_rd_en , 
    output reg  [6:0]  ram2_wr_addr, 
    output reg  [5:0]  ram2_rd_addr, 
    
    input  wire        data_en ,       
    input  wire [63:0] data_in ,       
    output reg         o_upstream_ready, 
    
    input  wire        i_downstream_ready, 
    output wire        o_data_valid,    
    output reg  [63:0] data_out            
);

    parameter   IDLE        = 4'b0001, 
                WRAM1       = 4'b0010, 
                WRAM2_RRAM1 = 4'b0100, 
                WRAM1_RRAM2 = 4'b1000; 

    // 写计数器�?大�?? 64
    localparam CNT_WR_MAX = 7'd64; 
    localparam CNT_RD_MAX = 6'd63; 

    reg [3:0] state ; 
    reg ram1_rd_done;
    reg ram2_rd_done;

    // ============================================================
    // 【关键修�?1】输入信号打�? (Register Input)
    // 解决 "data_in 不稳�?" 的问�?
    // ============================================================
    reg [63:0] data_in_d;
    reg        data_en_d;

    always @(posedge clk_50m or negedge rst_n) begin
        if(!rst_n) begin
            data_in_d <= 64'd0;
            data_en_d <= 1'b0;
        end
        else if(o_upstream_ready) begin
            // 只有�? Ready 为高时，才接收数据进寄存�?
            data_in_d <= data_in;
            data_en_d <= data_en;
        end
        else begin
            // 如果 Ready 拉低了，停止接收有效标志（防止溢出写入）
            data_en_d <= 1'b0;
        end
    end

    // ============================================================
    // 【关键修�?2】写数据使用打拍后的信号
    // ============================================================
    // 写数据源改为 data_in_d (寄存器输出，时序稳定)
    assign ram1_wr_data = (ram1_wr_en) ? data_in_d : 64'd0;
    assign ram2_wr_data = (ram2_wr_en) ? data_in_d : 64'd0;

    // ============================================================
    // 【关键修�?3】Ready 信号逻辑 (提前�?拍关�?)
    // ============================================================
    always @(*) begin
        case(state)
            IDLE:        o_upstream_ready = 1'b1; 
            
            // 注意：这里改成了 < 63 (CNT_WR_MAX - 1)
            // 为什么？因为我们加了寄存器延迟�??
            // �? ram_wr_addr 等于 63 时，说明 RAM 里已经写�? 63 个数�?
            // 但此时寄存器 data_in_d 里可能正存着�? 64 个数等待写入�?
            // �?以必须现在就拉低 Ready，阻止第 65 个数进入寄存器�??
            WRAM1:       o_upstream_ready = (ram1_wr_addr < (CNT_WR_MAX - 1'b1)); 
            WRAM1_RRAM2: o_upstream_ready = (ram1_wr_addr < (CNT_WR_MAX - 1'b1));
            WRAM2_RRAM1: o_upstream_ready = (ram2_wr_addr < (CNT_WR_MAX - 1'b1));
            
            default:     o_upstream_ready = 1'b0;
        endcase
    end

    // ============================================================
    // 写使能�?�辑 (使用打拍后的 Valid)
    // ============================================================
    always @(*) begin
        ram1_wr_en = 0;
        ram2_wr_en = 0;
        // 使用 data_en_d (延迟后的使能)
        // 注意：这里不�?要再判断 Ready，因�? data_en_d 的生成已经受 Ready 控制�?
        if(data_en_d) begin
            case(state)
                WRAM1, WRAM1_RRAM2: ram1_wr_en = 1;
                WRAM2_RRAM1:        ram2_wr_en = 1;
            endcase
        end
    end

    // ============================================================
    // 状�?�机 (保持 7 位计数器的跳转�?�辑)
    // ============================================================
    always@(posedge clk_50m or negedge rst_n)
        if(!rst_n) state <= IDLE;
        else case(state)
            IDLE: if(data_en) state <= WRAM1; // 这里可以�? data_en 或�?? data_en_d 启动，影响不�?
            
            // 只要地址到了 64，说明第 64 个数（存在寄存器里的那个）已经写进去�?
            WRAM1: if(ram1_wr_addr == CNT_WR_MAX) 
                       state <= WRAM2_RRAM1;
            
            WRAM2_RRAM1: if(ram2_wr_addr == CNT_WR_MAX && ram1_rd_done) 
                       state <= WRAM1_RRAM2;
            
            WRAM1_RRAM2: if(ram1_wr_addr == CNT_WR_MAX && ram2_rd_done) 
                       state <= WRAM2_RRAM1;
                       
            default: state <= IDLE;
        endcase

    // ============================================================
    // 写地�?逻辑 (7位计数器�?0~64)
    // ============================================================
    always@(posedge clk_50m or negedge rst_n) begin
        if(!rst_n) ram1_wr_addr <= 0;
        else if(state == WRAM2_RRAM1) ram1_wr_addr <= 0;
        else if(ram1_wr_en && ram1_wr_addr < CNT_WR_MAX) 
            ram1_wr_addr <= ram1_wr_addr + 1'b1;
    end

    always@(posedge clk_50m or negedge rst_n) begin
        if(!rst_n) ram2_wr_addr <= 0;
        else if(state == WRAM1_RRAM2 || state == WRAM1) ram2_wr_addr <= 0;
        else if(ram2_wr_en && ram2_wr_addr < CNT_WR_MAX) 
            ram2_wr_addr <= ram2_wr_addr + 1'b1;
    end

    // ============================================================
    // 读控制与输出 (保持原样)
    // ============================================================
    always @(*) begin
        ram1_rd_en = (state == WRAM2_RRAM1) && !ram1_rd_done;
        ram2_rd_en = (state == WRAM1_RRAM2) && !ram2_rd_done;
    end

    always@(posedge clk_50m or negedge rst_n) begin
        if(!rst_n) begin ram1_rd_addr <= 0; ram1_rd_done <= 0; end
        else if(state != WRAM2_RRAM1) begin ram1_rd_addr <= 0; ram1_rd_done <= 0; end
        else if(ram1_rd_en && i_downstream_ready) begin 
            if(ram1_rd_addr == CNT_RD_MAX) ram1_rd_done <= 1;
            else ram1_rd_addr <= ram1_rd_addr + 1'b1;
        end
    end

    always@(posedge clk_50m or negedge rst_n) begin
        if(!rst_n) begin ram2_rd_addr <= 0; ram2_rd_done <= 0; end
        else if(state != WRAM1_RRAM2) begin ram2_rd_addr <= 0; ram2_rd_done <= 0; end
        else if(ram2_rd_en && i_downstream_ready) begin 
            if(ram2_rd_addr == CNT_RD_MAX) ram2_rd_done <= 1;
            else ram2_rd_addr <= ram2_rd_addr + 1'b1;
        end
    end

    reg valid_reg;   
    always @(posedge clk_50m or negedge rst_n) begin
        if(!rst_n) 
            valid_reg <= 0;
        else if(i_downstream_ready)
            valid_reg <= (ram1_rd_en || ram2_rd_en);
    end
    assign o_data_valid = valid_reg && (ram1_rd_en || ram2_rd_en);

    always @(posedge clk_50m or negedge rst_n) begin
        if(!rst_n) 
            data_out <= 64'd0;
        else if(i_downstream_ready) begin
            if(ram1_rd_en)      data_out <= ram1_rd_data;
            else if(ram2_rd_en) data_out <= ram2_rd_data;
        end
    end

endmodule
//`timescale 1ns / 1ps
//module ram_ctrl1
//(
//    input  wire        clk_50m ,
//    input  wire        rst_n ,
    
//    input  wire [63:0] ram1_rd_data, 
//    input  wire [63:0] ram2_rd_data, 
//    output wire [63:0] ram1_wr_data, 
//    output wire [63:0] ram2_wr_data, 
    
//    output reg         ram1_wr_en , 
//    output reg         ram1_rd_en , 
    
//    output reg  [6:0]  ram1_wr_addr, 
//    output reg  [5:0]  ram1_rd_addr, 
    
//    output reg         ram2_wr_en , 
//    output reg         ram2_rd_en , 
//    output reg  [6:0]  ram2_wr_addr, 
//    output reg  [5:0]  ram2_rd_addr, 
    
//    input  wire        data_en ,       
//    input  wire [63:0] data_in ,     
//    input  wire        i_data_last,     // �������ݵĽ�����־  
//    output reg         o_upstream_ready, 
    
//    input  wire        i_downstream_ready, 
//    output wire        o_data_valid,    
//    output reg         o_data_last,     // ������ݵĽ�����־
//    output reg  [63:0] data_out            
//);

//    parameter   IDLE        = 4'b0001, 
//                WRAM1       = 4'b0010, 
//                WRAM2_RRAM1 = 4'b0100, 
//                WRAM1_RRAM2 = 4'b1000; 

//    localparam CNT_WR_MAX = 7'd64; 

//    reg [3:0] state ; 
//    reg ram1_rd_done;
//    reg ram2_rd_done;
    
//    // ��¼ÿ�� RAM ʵ��д������ݳ��� (1-64)
//    reg [6:0] ram1_len;
//    reg [6:0] ram2_len;

//    // ============================================================
//    // 1. �����źŴ���
//    // ============================================================
//    reg [63:0] data_in_d;
//    reg        data_en_d;
//    reg        i_data_last_d;

//    always @(posedge clk_50m or negedge rst_n) begin
//        if(!rst_n) begin
//            data_in_d <= 64'd0;
//            data_en_d <= 1'b0;
//            i_data_last_d <= 1'b0;
//        end
//        else if(o_upstream_ready) begin
//            data_in_d <= data_in;
//            data_en_d <= data_en;
//            i_data_last_d <= i_data_last;
//        end
//        else begin
//            data_en_d <= 1'b0;
//            i_data_last_d <= 1'b0;
//        end
//    end

//    assign ram1_wr_data = (ram1_wr_en) ? data_in_d : 64'd0;
//    assign ram2_wr_data = (ram2_wr_en) ? data_in_d : 64'd0;

//    // ============================================================
//    // 2. Ready �ź��߼� (��ǰһ�Ĺ���)
//    // ============================================================
//    always @(*) begin
//        case(state)
//            IDLE:        o_upstream_ready = 1'b1; 
//            WRAM1:       o_upstream_ready = (ram1_wr_addr < (CNT_WR_MAX - 1'b1)); 
//            WRAM1_RRAM2: o_upstream_ready = (ram1_wr_addr < (CNT_WR_MAX - 1'b1));
//            WRAM2_RRAM1: o_upstream_ready = (ram2_wr_addr < (CNT_WR_MAX - 1'b1));
//            default:     o_upstream_ready = 1'b0;
//        endcase
//    end

//    // ============================================================
//    // 3. ״̬�� (��������ж��볤�Ȳ���)
//    // ============================================================
//    always@(posedge clk_50m or negedge rst_n) begin
//        if(!rst_n) begin
//            state <= IDLE;
//            ram1_len <= 0;
//            ram2_len <= 0;
//        end
//        else case(state)
//            IDLE: if(data_en) state <= WRAM1; 
            
//            WRAM1: begin
//                // �����ַ�� 64 �����յ� last����ת����¼����
//                if(ram1_wr_en && (ram1_wr_addr == CNT_WR_MAX - 1'b1 || i_data_last_d)) begin
//                       state <= WRAM2_RRAM1;
//                       ram1_len <= ram1_wr_addr + 1'b1; 
//                end
//            end    

//            WRAM2_RRAM1: begin 
//                // ����������д��(���յ�last) �� ��һ�������Ѿ�����
//                if(ram2_wr_en && (ram2_wr_addr == CNT_WR_MAX - 1'b1 || i_data_last_d)) begin
//                    if(ram1_rd_done) begin // ���ֱ�������ֹ����δ������ RAM1
//                        state <= WRAM1_RRAM2;
//                        ram2_len <= ram2_wr_addr + 1'b1;
//                    end
//                end
//            end

//            WRAM1_RRAM2: begin 
//                if(ram1_wr_en && (ram1_wr_addr == CNT_WR_MAX - 1'b1 || i_data_last_d)) begin
//                    if(ram2_rd_done) begin // ���ֱ�������ֹ����δ������ RAM2
//                        state <= WRAM2_RRAM1;
//                        ram1_len <= ram1_wr_addr + 1'b1;
//                    end
//                end
//            end           
//            default: state <= IDLE;
//        endcase
//    end

//    // ============================================================
//    // 4. д��ַ�߼�
//    // ============================================================
//    always@(posedge clk_50m or negedge rst_n) begin
//        if(!rst_n) ram1_wr_addr <= 0;
//        else if(state == WRAM2_RRAM1) ram1_wr_addr <= 0;
//        else if(ram1_wr_en && ram1_wr_addr < CNT_WR_MAX) 
//            ram1_wr_addr <= ram1_wr_addr + 1'b1;
//    end

//    always@(posedge clk_50m or negedge rst_n) begin
//        if(!rst_n) ram2_wr_addr <= 0;
//        else if(state == WRAM1_RRAM2 || state == WRAM1) ram2_wr_addr <= 0;
//        else if(ram2_wr_en && ram2_wr_addr < CNT_WR_MAX) 
//            ram2_wr_addr <= ram2_wr_addr + 1'b1;
//    end

//    // ============================================================
//    // 5. �������߼� (��������ֹ�ж�)
//    // ============================================================
//    always @(*) begin
//        ram1_wr_en = (data_en_d && (state == WRAM1 || state == WRAM1_RRAM2));
//        ram2_wr_en = (data_en_d && (state == WRAM2_RRAM1));
//        ram1_rd_en = (state == WRAM2_RRAM1) && !ram1_rd_done;
//        ram2_rd_en = (state == WRAM1_RRAM2) && !ram2_rd_done;
//    end

//    always@(posedge clk_50m or negedge rst_n) begin
//        if(!rst_n) begin ram1_rd_addr <= 0; ram1_rd_done <= 0; end
//        else if(state != WRAM2_RRAM1) begin ram1_rd_addr <= 0; ram1_rd_done <= 0; end
//        else if(ram1_rd_en && i_downstream_ready) begin 
//            // �������Ա�ʵ�ʳ��� ram1_len������������ 63
//            if(ram1_rd_addr == ram1_len[5:0] - 1'b1) 
//                ram1_rd_done <= 1;
//            else 
//                ram1_rd_addr <= ram1_rd_addr + 1'b1;
//        end
//    end

//    always@(posedge clk_50m or negedge rst_n) begin
//        if(!rst_n) begin ram2_rd_addr <= 0; ram2_rd_done <= 0; end
//        else if(state != WRAM1_RRAM2) begin ram2_rd_addr <= 0; ram2_rd_done <= 0; end
//        else if(ram2_rd_en && i_downstream_ready) begin 
//            if(ram2_rd_addr == ram2_len[5:0] - 1'b1) 
//                ram2_rd_done <= 1;
//            else 
//                ram2_rd_addr <= ram2_rd_addr + 1'b1;
//        end
//    end

//    // ============================================================
//    // 6. ��� Valid/Last/Data (���߶���)
//    // ============================================================
//    reg valid_reg;   
//    always @(posedge clk_50m or negedge rst_n) begin
//        if(!rst_n) begin
//            valid_reg <= 0;
//            o_data_last <= 0;
//        end
//        else if(i_downstream_ready) begin
//            valid_reg   <= (ram1_rd_en || ram2_rd_en);
//            // Last �� Valid ͬ�����Ĳ���
//            o_data_last <= (ram1_rd_en && (ram1_rd_addr == ram1_len[5:0] - 1'b1)) || 
//                           (ram2_rd_en && (ram2_rd_addr == ram2_len[5:0] - 1'b1));
//        end
//    end
//    assign o_data_valid = valid_reg;

//    always @(posedge clk_50m or negedge rst_n) begin
//        if(!rst_n) 
//            data_out <= 64'd0;
//        else if(i_downstream_ready) begin
//            if(ram1_rd_en)      data_out <= ram1_rd_data;
//            else if(ram2_rd_en) data_out <= ram2_rd_data;
//        end
//    end

//endmodule