`timescale 1ns / 1ps

module system_top(
    input  wire        sys_clk,
    input  wire        sys_rst_n,
    
    // === �ⲿ���� (ģ�� DMA) ===
    input  wire        dma_valid,      // Valid
    input  wire [63:0] dma_data,       // Data
    output wire        dma_ready,      // Ready (��ѹ����� DMA)
   // ===  ��̬���ýӿ� (����) === 
    input  wire [15:0] cfg_width,    // ���� 224
    input  wire [15:0] cfg_height,   // ���� 224
    input  wire        cfg_pad_en,
    // === �ⲿ��� (ģ�� ����˽ӿ�) ===
    output wire        conv_valid,     
    output wire [575:0] conv_window    // 3x3 * 8ch * 8bit
);

    // --- �ڲ������ź� ---
    wire [63:0] pp_data_out;    
    wire        pp_valid_out;   
    wire        padding_ready;  // ���ؼ�����������ź��� Padding ��������

    // ============================================================
    // 1. ʵ���� Ping-Pong Buffer (���뻺��)
    // ============================================================
    pingpang u_pingpang (
        .sys_clk            (sys_clk),
        .sys_rst_n          (sys_rst_n),
        
        // ���νӿ� (DMA <-> PingPang)
        .data_en            (dma_valid),
        .data_in            (dma_data),
        .o_upstream_ready   (dma_ready),
        
        // ���νӿ� (PingPang <-> Padding)
        .i_downstream_ready (padding_ready), // �������� Padding �ķ�ѹ
        .o_downstream_valid (pp_valid_out),
        .data_out           (pp_data_out)
    );

    // ============================================================
    // 2. ʵ���� Padding Module (��������)
    // ============================================================
    // �������Ѿ��� padding.v ������� output wire o_ready
    
    padding #(
        .NUM_CHANNELS (8),
        .DATA_WIDTH   (8),
        .MAX_IMG_WIDTH(1024),
        .FILTER_SIZE  (3)
    ) u_padding (
        .clk             (sys_clk),
        .rst_n           (sys_rst_n),
        // ������        
        .i_cfg_width     (cfg_width),
        .i_cfg_height    (cfg_height),
        .i_cfg_pad_en    (cfg_pad_en     ),
        .i_valid         (pp_valid_out),
        .i_data_parallel (pp_data_out),
        .o_ready         (padding_ready), // ���ؼ������ӷ�ѹ���
        
        // �����
        .o_valid         (conv_valid),
        .o_windows_packed(conv_window)
    );

endmodule
