`timescale 1ns / 1ps

module tb_line_buffer_with_padding;

    // =================================================================
    // 1. ����������� (��С�ߴ��Ա�۲�)
    // =================================================================
    parameter NUM_CHANNELS = 2;   // ����2��ͨ�������ڹ۲�
    parameter DATA_WIDTH   = 8;
    parameter IMG_WIDTH    = 5;   // 5x5 ��Сͼ
    parameter IMG_HEIGHT   = 5;
    parameter FILTER_SIZE  = 3;
    
    // =================================================================
    // 2. �źŶ���
    // =================================================================
    reg clk;
    reg rst_n;
    reg i_valid;
    reg [NUM_CHANNELS*DATA_WIDTH-1:0] i_data_parallel;
    
    wire o_valid;
    wire [NUM_CHANNELS*FILTER_SIZE*FILTER_SIZE*DATA_WIDTH-1:0] o_windows_packed;

    // =================================================================
    // 3. ����ģ��ʵ���� (DUT)
    // =================================================================
    line_buffer_with_padding #(
        .NUM_CHANNELS (NUM_CHANNELS),
        .DATA_WIDTH   (DATA_WIDTH),
        .IMG_WIDTH    (IMG_WIDTH),
        .IMG_HEIGHT   (IMG_HEIGHT),
        .FILTER_SIZE  (FILTER_SIZE)
    ) dut (
        .clk              (clk),
        .rst_n            (rst_n),
        .i_valid          (i_valid),
        .i_data_parallel  (i_data_parallel),
        .o_valid          (o_valid),
        .o_windows_packed (o_windows_packed)
    );

    // =================================================================
    // 4. ʱ������
    // =================================================================
    initial begin
        clk = 0;
        forever #5 clk = ~clk; // 10ns ����
    end

    // =================================================================
    // 5. ���Լ��� (Stimulus)
    // =================================================================
    integer r, c, ch;
    
    // �������ɲ�������ֵ�ĸ��������� Channel 0 = row*10 + col, Channel 1 = 0xFF
    function [DATA_WIDTH-1:0] get_pixel_val(input integer row, input integer col, input integer chan);
        if (chan == 0)
            get_pixel_val = (row * 10) + col; // ͨ��0��ֱ�۵�����ֵ (���� 12 �����1�е�2��)
        else
            get_pixel_val = 8'hFF;            // ͨ��1��ȫ1����������
    endfunction

    initial begin
        // --- ��ʼ�� ---
        rst_n = 0;
        i_valid = 0;
        i_data_parallel = 0;
        
        // --- �������μ�¼ (���ʹ�� Vivado/ModelSim) ---
        $dumpfile("wave.vcd");
        $dumpvars(0, tb_line_buffer_with_padding);

        // --- ��λ�ͷ� ---
        #20;
        rst_n = 1;
        #10;

        $display("-------------------------------------------------------------");
        $display("Simulation Start: Image Size %0dx%0d", IMG_WIDTH, IMG_HEIGHT);
        $display("-------------------------------------------------------------");

        // --- �������з������� ---
        // Ϊ��ȷ����ˮ����ȫ��������ǿ�����Ҫ�෢��һЩ��Ч���ڻ�Flush��
        // ����������߼���ֻҪʱ�����ܣ��л���ͻ�������
        // ���������ϸ��� 5x5 �������ݡ�
        
        for (r = 0; r < IMG_HEIGHT; r = r + 1) begin
            for (c = 0; c < IMG_WIDTH; c = c + 1) begin
                
                // �����ͨ����������
                for (ch = 0; ch < NUM_CHANNELS; ch = ch + 1) begin
                    i_data_parallel[ch*DATA_WIDTH +: DATA_WIDTH] = get_pixel_val(r, c, ch);
                end
                
                i_valid = 1;
                
                // ��ӡ������־
                if (ch == 0) // ����ӡ������Ϣ����ˢ��
                    $display("Input  @ Time %0t: Row=%0d, Col=%0d, Val_Ch0=%02d", $time, r, c, get_pixel_val(r,c,0));
                
                #10; // �ȴ�һ��ʱ������
            end
        end

        // --- �������룬��������ʱ���Թ۲�ʣ����� ---
        i_valid = 0;
        i_data_parallel = 0;
        
        #200; // �ȴ��㹻��ʱ������ˮ���ſ� (Padding Bottom��Ҫʱ��)
        
        $display("-------------------------------------------------------------");
        $display("Simulation Done");
        $finish;
    end

    // =================================================================
    // 6. ������ (Monitor)
    // =================================================================
    // ���� Packed �����Ա��ӡ
    reg [DATA_WIDTH-1:0] debug_window [NUM_CHANNELS-1:0][FILTER_SIZE-1:0][FILTER_SIZE-1:0];
    
    integer i, j, k;
    always @(*) begin
        for (i = 0; i < NUM_CHANNELS; i = i + 1) begin
            for (j = 0; j < FILTER_SIZE; j = j + 1) begin
                for (k = 0; k < FILTER_SIZE; k = k + 1) begin
                    debug_window[i][j][k] = o_windows_packed[ (i*9 + j*3 + k)*DATA_WIDTH +: DATA_WIDTH ];
                end
            end
        end
    end

    // ֻ�е� valid ��Чʱ�Ŵ�ӡ��������
    always @(posedge clk) begin
        if (o_valid) begin
            $display(">> OUTPUT VALID @ Time %0t", $time);
            // ��ӡ Channel 0 �� 3x3 ����
            $display("   [Channel 0 Window]:");
            $display("   %2d %2d %2d", debug_window[0][0][0], debug_window[0][0][1], debug_window[0][0][2]);
            $display("   %2d %2d %2d", debug_window[0][1][0], debug_window[0][1][1], debug_window[0][1][2]);
            $display("   %2d %2d %2d", debug_window[0][2][0], debug_window[0][2][1], debug_window[0][2][2]);
            $display("");
        end
    end

endmodule

