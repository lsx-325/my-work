// `timescale 1ns / 1ps

// module padding #(
//     parameter NUM_CHANNELS = 8,    
//     parameter DATA_WIDTH   = 64,    
//     parameter IMG_WIDTH    = 512,    
//     parameter IMG_HEIGHT   = 512,    
//     parameter FILTER_SIZE  = 3     
// )(
//     input                                   clk,
//     input                                   rst_n,
//     input                                   i_cfg_pad_en, // 1=����Padding(Same), 0=�ر�(Valid)
//     input                                   i_valid,
//     input [NUM_CHANNELS*DATA_WIDTH-1:0]     i_data_parallel,

//     output reg                              o_valid,
//     output wire                             o_ready, // ���������������Σ��ҿ��Խ�������
//     output [NUM_CHANNELS*FILTER_SIZE*FILTER_SIZE*DATA_WIDTH-1:0] o_windows_packed
// );

//     // 1. ��������
//     localparam PAD = FILTER_SIZE / 2; 
//     localparam TOTAL_WIDTH  = IMG_WIDTH + 2*PAD; 
//     localparam TOTAL_HEIGHT = IMG_HEIGHT + 2*PAD; 

//     // 2. FWFT FIFO
//     wire [NUM_CHANNELS*DATA_WIDTH-1:0] fifo_dout;
//     wire fifo_empty;
//     reg  fifo_rd_en;
//     wire fifo_full;
    
//     fwft_fifo_behavioral #(.DATA_WIDTH(NUM_CHANNELS*DATA_WIDTH), .DEPTH(512)) u_input_fifo (
//         .clk(clk), .rst_n(rst_n),
//         .wr_en(i_valid), .din(i_data_parallel),
//         .rd_en(fifo_rd_en), .dout(fifo_dout),
//         .empty(fifo_empty), .full(fifo_full)
//     );
//     assign o_ready = !fifo_full; // ����� Ping-Pong

//     // 3. ɨ��״̬��
//     reg [15:0] x_cnt, y_cnt; 
//     reg running; 
//     wire in_active_region = (x_cnt >= PAD) && (x_cnt < IMG_WIDTH + PAD) && (y_cnt >= PAD) && (y_cnt < IMG_HEIGHT + PAD);
//     wire can_advance = in_active_region ? (!fifo_empty) : 1'b1;

//     always @(*) fifo_rd_en = (in_active_region && !fifo_empty) ? 1'b1 : 1'b0;

//     always @(posedge clk or negedge rst_n) begin
//         if (!rst_n) begin
//             x_cnt <= 0; y_cnt <= 0; running <= 0;
//         end else begin
//             if (!fifo_empty) running <= 1; 
//             if (running && can_advance) begin
//                 if (x_cnt == TOTAL_WIDTH - 1) begin
//                     x_cnt <= 0;
//                     if (y_cnt == TOTAL_HEIGHT - 1) begin y_cnt <= 0; running <= 0; end 
//                     else y_cnt <= y_cnt + 1;
//                 end else x_cnt <= x_cnt + 1;
//             end
//         end
//     end

//     // 4. ������ (������ˮ�� d2����֤��ֱ����)
//     reg [NUM_CHANNELS*DATA_WIDTH-1:0] current_stream_pixel;
//     reg [NUM_CHANNELS*DATA_WIDTH-1:0] current_stream_pixel_d1; 
//     reg [NUM_CHANNELS*DATA_WIDTH-1:0] current_stream_pixel_d2; 
//     reg                               current_stream_valid;

//     always @(posedge clk or negedge rst_n) begin
//         if (!rst_n) begin
//             current_stream_pixel <= 0; 
//             current_stream_pixel_d1 <= 0; 
//             current_stream_pixel_d2 <= 0;
//             current_stream_valid <= 0;
//         end else if (running && can_advance) begin
//             current_stream_valid <= 1;
//             // Stage 0
//             if (in_active_region) current_stream_pixel <= fifo_dout; else current_stream_pixel <= 0;
//             // Stage 1
//             current_stream_pixel_d1 <= (in_active_region) ? fifo_dout : 0;
//             // Stage 2 (Window Input)
//             current_stream_pixel_d2 <= current_stream_pixel_d1;
//         end else begin
//             current_stream_valid <= 0;
//         end
//     end

//     // 5. Line Buffers
//     reg [NUM_CHANNELS*DATA_WIDTH-1:0] lb0 [0:TOTAL_WIDTH-1]; 
//     reg [NUM_CHANNELS*DATA_WIDTH-1:0] lb1 [0:TOTAL_WIDTH-1]; 
//     reg [NUM_CHANNELS*DATA_WIDTH-1:0] rdata_lb0, rdata_lb1;
//     reg [15:0] x_cnt_d1;
//     integer i;
//     initial begin for (i=0; i<TOTAL_WIDTH; i=i+1) begin lb0[i] = 0; lb1[i] = 0; end end

//     always @(posedge clk or negedge rst_n) begin
//         if (!rst_n) begin
//             rdata_lb0 <= 0; rdata_lb1 <= 0; x_cnt_d1 <= 0;
//             for (i=0; i<TOTAL_WIDTH; i=i+1) begin lb0[i] <= 0; lb1[i] <= 0; end
//         end else if (running && can_advance) begin
//             x_cnt_d1 <= x_cnt;
//             rdata_lb0 <= lb0[x_cnt]; rdata_lb1 <= lb1[x_cnt];
//             lb0[x_cnt] <= current_stream_pixel; lb1[x_cnt_d1] <= rdata_lb0; 
//         end
//     end

//     // 6. ���� & ���� Valid ����
//     reg [NUM_CHANNELS*DATA_WIDTH-1:0] win [0:2][0:2]; 
//     integer r, c;
    
//     reg ramp_up_done;
//     always @(posedge clk or negedge rst_n) begin
//         if(!rst_n) ramp_up_done <= 0;
//         else if (y_cnt == 2) ramp_up_done <= 1; 
//         else if (!running) ramp_up_done <= 0;
//     end

//     // === ������� Valid �ж� (������� 1 ��) ===
    
//     // Phase A: ɨ���е�ǰ��� (x=4, 5) -> ��Ӧ Pixel 1, 2
//     wire phase_a_x = (x_cnt == 4 || x_cnt == 5);
//     wire phase_a_y = (y_cnt >= 2 && y_cnt <= 5);

//     // Phase B: ɨ���еĺ��� (x=0, 1) -> ��Ӧ Pixel 3, 4
//     // ע�⣺�޳��� x=2 (Right Pad)
//     wire phase_b_x = (x_cnt == 0 || x_cnt == 1);
//     wire phase_b_y = (y_cnt >= 3 || y_cnt == 0);

//     always @(posedge clk or negedge rst_n) begin
//         if (!rst_n) begin
//             o_valid <= 0;
//             for(r=0; r<3; r=r+1) for(c=0; c<3; c=c+1) win[r][c] <= 0;
//         end else if (current_stream_valid) begin
//             for(r=0; r<3; r=r+1) for(c=0; c<2; c=c+1) win[r][c] <= win[r][c+1];
            
//             win[2][2] <= current_stream_pixel_d2; 
//             win[1][2] <= rdata_lb0; 
//             win[0][2] <= rdata_lb1;

//             if ( ramp_up_done && ( (phase_a_x && phase_a_y) || (phase_b_x && phase_b_y) ) ) 
//                 o_valid <= 1;
//             else
//                 o_valid <= 0;
//         end else begin
//             o_valid <= 0;
//         end
//     end

//     // 7. ��� (����)
//     genvar gr, gc;
//     generate
//         for (gr = 0; gr < 3; gr = gr + 1) begin : pack_row
//             for (gc = 0; gc < 3; gc = gc + 1) begin : pack_col
//                 assign o_windows_packed[((gr*3 + gc + 1)*NUM_CHANNELS*DATA_WIDTH)-1 -: NUM_CHANNELS*DATA_WIDTH] 
//                        = win[gr][gc];
//             end
//         end
//     endgenerate
// endmodule

// // FWFT FIFO Module (Same as before)
// module fwft_fifo_behavioral #(
//     parameter DATA_WIDTH = 64, 
//     parameter DEPTH = 512)(
//     input clk, rst_n, wr_en, 
//     input [DATA_WIDTH-1:0] din, 
//     input rd_en,
//     output [DATA_WIDTH-1:0] dout, 
//     output empty, 
//     output full
// );
//     reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];
//     reg [15:0] wr_ptr = 0, rd_ptr = 0, count = 0;
//     assign empty = (count == 0); assign full  = (count == DEPTH);
//     assign dout = mem[rd_ptr];
//     always @(posedge clk or negedge rst_n) begin
//         if (!rst_n) begin wr_ptr<=0; rd_ptr<=0; count<=0; end
//         else begin
//             if (wr_en && !full) begin
//                 mem[wr_ptr] <= din; wr_ptr <= (wr_ptr==DEPTH-1)?0:wr_ptr+1;
//                 if (!rd_en) count <= count + 1;
//             end
//             if (rd_en && !empty) begin
//                 rd_ptr <= (rd_ptr==DEPTH-1)?0:rd_ptr+1;
//                 if (!wr_en) count <= count - 1;
//             end
//         end
//     end
// endmodule
`timescale 1ns / 1ps

module padding #(
    parameter NUM_CHANNELS = 8,    
    parameter DATA_WIDTH   = 8,    
    // ��Ӳ����Դ���ޡ����� >= ʵ���������
    parameter MAX_IMG_WIDTH = 1024, 
    parameter FILTER_SIZE  = 3     
)(
    input                                   clk,
    input                                   rst_n,
    
    // === ��̬���ýӿ� ===
    input [15:0]                            i_cfg_width ,  // ��ǰ��� (e.g. 4, 224, 512)
    input [15:0]                            i_cfg_height, // ��ǰ���
    input                                   i_cfg_pad_en, // 1=����Padding(Same), 0=�ر�(Valid)
    
    // === �������ӿ� ===
    input                                   i_valid,
    input [NUM_CHANNELS*DATA_WIDTH-1:0]     i_data_parallel,
    output reg                              o_valid,
    output wire                             o_ready,      // ��ѹ�ź�
    output [NUM_CHANNELS*FILTER_SIZE*FILTER_SIZE*DATA_WIDTH-1:0] o_windows_packed
);

    // ============================================================
    // 1. �����밲ȫ����
    // ============================================================
    localparam PAD = FILTER_SIZE / 2; 

    // ����ȫ�������������ÿ�Ȳ�����Ӳ�����ޣ���ֹ BRAM ���
    wire [15:0] safe_cfg_width = (i_cfg_width > MAX_IMG_WIDTH) ? MAX_IMG_WIDTH : i_cfg_width;

    // ��̬�����ܳߴ� (Image + Padding)
    wire [15:0] total_width  = safe_cfg_width + 2*PAD; 
    wire [15:0] total_height = i_cfg_height + 2*PAD; 

    // ============================================================
    // 2. ���뻺�� FIFO (FWFT)
    // ============================================================
    wire [NUM_CHANNELS*DATA_WIDTH-1:0] fifo_dout;
    wire fifo_empty, fifo_full;
    reg  fifo_rd_en;

    fwft_fifo_behavioral #(.DATA_WIDTH(NUM_CHANNELS*DATA_WIDTH), .DEPTH(1024)) u_input_fifo (
        .clk(clk), .rst_n(rst_n),
        .wr_en(i_valid), .din(i_data_parallel),
        .rd_en(fifo_rd_en), .dout(fifo_dout),
        .empty(fifo_empty), .full(fifo_full)
    );
    // �����ѹ�ź�
    assign o_ready = !fifo_full; 

    // ============================================================
    // 3. ����ɨ��״̬��
    // ============================================================
    reg [15:0] x_cnt, y_cnt; 
    reg running; 
    
    // �жϵ�ǰɨ����Ƿ���"��Чͼ������"�� (���ھ����Ǵ� FIFO �����ݻ��ǲ� 0)
    wire in_active_region = (x_cnt >= PAD) && (x_cnt < safe_cfg_width + PAD) && 
                            (y_cnt >= PAD) && (y_cnt < i_cfg_height + PAD);
                            
    // ֻҪ������Ч�����ڣ�����Ҫ FIFO �����ݲ���ǰ��������(��Padding��)����ֱ����
    wire can_advance = in_active_region ? (!fifo_empty) : 1'b1;

    always @(*) fifo_rd_en = (in_active_region && !fifo_empty) ? 1'b1 : 1'b0;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            x_cnt <= 0; y_cnt <= 0; running <= 0;
        end else begin
            if (!fifo_empty) running <= 1; 
            if (running && can_advance) begin
                // ���� Total Width ɨ��
                if (x_cnt == total_width - 1) begin
                    x_cnt <= 0;
                    if (y_cnt == total_height - 1) begin y_cnt <= 0; running <= 0; end 
                    else y_cnt <= y_cnt + 1;
                end else x_cnt <= x_cnt + 1;
            end
        end
    end

    // ============================================================
    // 4. �л��� (Line Buffers)
    // ============================================================
    reg [NUM_CHANNELS*DATA_WIDTH-1:0] current_stream_pixel;
    reg [NUM_CHANNELS*DATA_WIDTH-1:0] current_stream_pixel_d2; 
    reg                               current_stream_valid;

    // BRAM ��Դ����
    localparam LB_DEPTH = MAX_IMG_WIDTH + 2*PAD; 
    reg [NUM_CHANNELS*DATA_WIDTH-1:0] lb0 [0:LB_DEPTH-1]; 
    reg [NUM_CHANNELS*DATA_WIDTH-1:0] lb1 [0:LB_DEPTH-1]; 
    reg [NUM_CHANNELS*DATA_WIDTH-1:0] rdata_lb0, rdata_lb1;

    always @(posedge clk) begin
        if (running && can_advance) begin
            // 1. �ȶ�����ǰλ�õľ����� (���ڻ������м��кͶ���)
            rdata_lb0 <= lb0[x_cnt];
            rdata_lb1 <= lb1[x_cnt];
            
            // 2. ׼�������� (���� FIFO �� Padding 0)
            if (in_active_region) current_stream_pixel <= fifo_dout; 
            else current_stream_pixel <= 0;

            // 3. д�� Line Buffer (���»���)
            // LB0 �������У�LB1 �������(�� rdata_lb0)
            lb0[x_cnt] <= (in_active_region) ? fifo_dout : 0; 
            // ע�⣺�������ǰ���һ�Ĵ��� lb0 ������(���ڶ������� rdata_lb0) ���� lb1
            // ������ʱ���߼�����ͬһ��ʹ�� lb0[x_cnt] (����ǰ) ����ֱ�ӵ���λ��ʽ
            lb1[x_cnt] <= lb0[x_cnt]; 
        end
    end

    // ������ˮ���ӳ� (Input -> Window Bottom ��Ҫƥ�� RAM ��ȡ�ӳ�)
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin 
            current_stream_valid <= 0; 
            current_stream_pixel_d2 <= 0;
        end else if (running && can_advance) begin
            current_stream_valid <= 1;
            current_stream_pixel_d2 <= (in_active_region) ? fifo_dout : 0; 
        end else begin
            current_stream_valid <= 0;
        end
    end

    // ============================================================
    // 5. �������ڹ��� (3x3 Shift Register)
    // ============================================================
    reg [NUM_CHANNELS*DATA_WIDTH-1:0] win [0:2][0:2]; 
    integer r, c;
    reg ramp_up_done;
    
    // Ԥ���߼����ȴ�ǰ�����������ҵ����е�ǰ�������ؽ�����λ�Ĵ���
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) ramp_up_done <= 0;
        else if (y_cnt == 2 && x_cnt == 2) ramp_up_done <= 1; 
        else if (!running) ramp_up_done <= 0;
    end
    
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
             for(r=0; r<3; r=r+1) for(c=0; c<3; c=c+1) win[r][c] <= 0;
        end else if (current_stream_valid) begin
             // ���Ʋ���
             for(r=0; r<3; r=r+1) for(c=0; c<2; c=c+1) win[r][c] <= win[r][c+1];
             // �µ�һ�н���
             win[2][2] <= current_stream_pixel_d2; // Bottom
             win[1][2] <= rdata_lb0;                 // Middle
             win[0][2] <= rdata_lb1;                 // Top
        end
    end

    // ============================================================
    // 6. [������] �������׷���� Valid �ж�
    // ============================================================
    reg [15:0] out_x, out_y;

    // 6.1 ���������
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            out_x <= 0; out_y <= 0; 
        end else if (current_stream_valid && ramp_up_done) begin
            // ���� Total Width ѭ������
            if (out_x == total_width - 1) begin
                out_x <= 0;
                if (out_y == total_height - 1) out_y <= 0;
                else out_y <= out_y + 1;
            end else begin
                out_x <= out_x + 1;
            end
        end else if (!running) begin
             out_x <= 0; out_y <= 0;
        end
    end

    // 6.2 ��Ե����Ч���ж� (��Ϊ����߼� Wire������1���ӳ٣����Center=1��ʧ����)
    
    // �жϵ�ǰ���Ƿ�������Чͼ������ (0 ~ width-1)
    wire is_active_col = (out_x < safe_cfg_width); 
    
    // ��Ե�ж�
    wire is_border_left   = (out_x == 0);
    wire is_border_right  = (out_x == safe_cfg_width - 1);
    wire is_border_top    = (out_y == 0);
    wire is_border_bottom = (out_y == i_cfg_height - 1);
    wire is_border = is_border_left || is_border_right || is_border_top || is_border_bottom;

    // 6.3 ������� Valid ����
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            o_valid <= 0;
        end else if (current_stream_valid && ramp_up_done) begin
            // ֻ�е���ǰ������Чͼ������ʱ���ſ������ Valid
            // (���˵���βΪ�˲��� Padding ����������������)
            if (is_active_col) begin
                if (i_cfg_pad_en) begin
                    // ������ Padding��: ���������Ч�У�������Ե
                    o_valid <= 1'b1;
                end else begin
                    // ���ر� Padding��: ����Ǳ�Ե������
                    if (is_border) 
                        o_valid <= 1'b0;
                    else 
                        o_valid <= 1'b1;
                end
            end else begin
                o_valid <= 1'b0;
            end
        end else begin
            o_valid <= 0;
        end
    end

    // ============================================================
    // 7. ������
    // ============================================================
    genvar gr, gc;
    generate
        for (gr = 0; gr < 3; gr = gr + 1) begin : pack_row
            for (gc = 0; gc < 3; gc = gc + 1) begin : pack_col
                assign o_windows_packed[((gr*3 + gc + 1)*NUM_CHANNELS*DATA_WIDTH)-1 -: NUM_CHANNELS*DATA_WIDTH] 
                       = win[gr][gc];
            end
        end
    endgenerate

endmodule

// ============================================================
// ����FWFT FIFO ģ�� (�������)
// ============================================================
module fwft_fifo_behavioral #(
    parameter DATA_WIDTH = 64, 
    parameter DEPTH = 512)(
    input clk, rst_n, wr_en, 
    input [DATA_WIDTH-1:0] din, 
    input rd_en,
    output [DATA_WIDTH-1:0] dout, 
    output empty, 
    output full
);
    reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];
    reg [15:0] wr_ptr = 0, rd_ptr = 0, count = 0;
    
    assign empty = (count == 0); 
    assign full  = (count == DEPTH);
    assign dout = mem[rd_ptr]; // FWFT ���ԣ�����ֱ�����
    
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin wr_ptr<=0; rd_ptr<=0; count<=0; end
        else begin
            if (wr_en && !full) begin
                mem[wr_ptr] <= din; 
                wr_ptr <= (wr_ptr==DEPTH-1)?0:wr_ptr+1;
                if (!rd_en) count <= count + 1;
            end
            if (rd_en && !empty) begin
                rd_ptr <= (rd_ptr==DEPTH-1)?0:rd_ptr+1;
                if (!wr_en) count <= count - 1;
            end
        end
    end
endmodule