//`timescale 1ns / 1ps

//module tb_fpga_top_level_new;

//    // =========================================================================
//    // 1. ��������
//    // =========================================================================
//    parameter AXIS_DATA_WIDTH = 64;
//    parameter NUM_IN_CHANNELS = 8;
//    parameter DATA_WIDTH      = 8;
//    parameter ACCUM_WIDTH     = 32;
//    parameter FILTER_SIZE     = 3;
    
//    // Ϊ�˷����ٶȣ����ǽ�ͼ��ߴ���Сһ��
//    parameter IMG_WIDTH       = 16; 
//    parameter IMG_HEIGHT      = 16;
//    parameter BRAM_DEPTH      = 512;

//    // Ȩ�ؼ�����ؼ���
//    // Layer 1: 4 Cores, ÿ�� Core ���� 2 �����ͨ��
//    // ÿ�� Core ��Ҫ 144 ��Ȩ�� (8 In * 2 Out * 9) = 1152 bits
//    // 1152 bits / 64 bits (AXI) = 18 Beats
//    parameter BEATS_PER_WEIGHT_LINE = (NUM_IN_CHANNELS * 2 * FILTER_SIZE * FILTER_SIZE * DATA_WIDTH) / AXIS_DATA_WIDTH;

//    // =========================================================================
//    // 2. �źŶ���
//    // =========================================================================
//    reg clk;
//    reg rst_n;

//    // ͼ������
//    reg                       s_axis_img_tvalid;
//    wire                      s_axis_img_tready;
//    reg [AXIS_DATA_WIDTH-1:0] s_axis_img_tdata;
//    reg                       s_axis_img_tlast;

//    // Ȩ������
//    reg                       s_axis_w_tvalid;
//    wire                      s_axis_w_tready;
//    reg [AXIS_DATA_WIDTH-1:0] s_axis_w_tdata;
//    reg                       s_axis_w_tlast;

//    // ������
//    wire                      m_axis_res_tvalid;
//    reg                       m_axis_res_tready;
//    wire [AXIS_DATA_WIDTH-1:0] m_axis_res_tdata;
//    wire [AXIS_DATA_WIDTH/8-1:0] m_axis_res_tkeep;
//    wire                      m_axis_res_tlast;

//    // �����ź�
//    reg                       i_load_weights;
//    reg [3:0]                 i_target_layer;
//    reg                       i_start_compute;
//    reg [8:0]                 i_l1_weight_base;
//    reg [8:0]                 i_l2_weight_base;
//    wire                      o_compute_done;

//    // ͳ�ƽ��յ���������
//    integer received_pixel_cnt;
//    integer k, r, c, pixel_idx;

//    // =========================================================================
//    // 3. DUT ʵ����
//    // =========================================================================
//    fpga_top_level #(
//        .AXIS_DATA_WIDTH(AXIS_DATA_WIDTH),
//        .NUM_IN_CHANNELS(NUM_IN_CHANNELS),
//        .DATA_WIDTH     (DATA_WIDTH),
//        .ACCUM_WIDTH    (ACCUM_WIDTH),
//        .FILTER_SIZE    (FILTER_SIZE),
//        .IMG_WIDTH      (IMG_WIDTH),
//        .IMG_HEIGHT     (IMG_HEIGHT),
//        .BRAM_DEPTH     (BRAM_DEPTH)
//    ) u_dut (
//        .clk(clk),
//        .rst_n(rst_n),
        
//        .s_axis_img_tvalid(s_axis_img_tvalid),
//        .s_axis_img_tready(s_axis_img_tready),
//        .s_axis_img_tdata (s_axis_img_tdata),
//        .s_axis_img_tlast (s_axis_img_tlast),
        
//        .s_axis_w_tvalid  (s_axis_w_tvalid),
//        .s_axis_w_tready  (s_axis_w_tready),
//        .s_axis_w_tdata   (s_axis_w_tdata),
//        .s_axis_w_tlast   (s_axis_w_tlast),
        
//        .m_axis_res_tvalid(m_axis_res_tvalid),
//        .m_axis_res_tready(m_axis_res_tready),
//        .m_axis_res_tdata (m_axis_res_tdata),
//        .m_axis_res_tkeep (m_axis_res_tkeep),
//        .m_axis_res_tlast (m_axis_res_tlast),
        
//        .i_load_weights   (i_load_weights),
//        .i_target_layer   (i_target_layer),
//        .i_start_compute  (i_start_compute),
//        .i_l1_weight_base (i_l1_weight_base),
//        .i_l2_weight_base (i_l2_weight_base),
//        .o_compute_done   (o_compute_done)
//    );

//    // =========================================================================
//    // 4. ʱ������ (100MHz)
//    // =========================================================================
//    initial begin
//        clk = 0;
//        forever #5 clk = ~clk;
//    end

//    // =========================================================================
//    // 5. ������ (Helper Tasks)
//    // =========================================================================
    
//    // ���񣺼���һ��Ȩ�ص�ָ���� Target Layer
//    task load_weights_for_target;
//        input [3:0] target_id;
//        input [7:0] start_val;
        
//        reg [7:0] k_val;
//        begin
//            $display("[Time %0t] Loading Weights for Target ID: %d", $time, target_id);
            
//            // 1. ���ÿ����ź�
//            @(posedge clk);
//            i_target_layer = target_id;
//            i_load_weights = 1; // ������λ����
//            @(posedge clk);
//            i_load_weights = 0; // �������壬��ʼ����
            
//            // 2. ���� AXI Stream ����
//            // ����ÿ�� Core ֻ��Ҫ 1 ��Ȩ�� (Addr 0)����Ҫ���� BEATS_PER_WEIGHT_LINE ��
//            for (k = 0; k < BEATS_PER_WEIGHT_LINE; k = k + 1) begin
//                s_axis_w_tvalid = 1;
//                k_val = start_val + k;
//                // ����������ݣ��򵥵ĵ��������������
//                s_axis_w_tdata  = {8{k_val}}; 
                
//                if (k == BEATS_PER_WEIGHT_LINE - 1) 
//                    s_axis_w_tlast = 1;
//                else 
//                    s_axis_w_tlast = 0;
                
//                @(posedge clk);
//            end
            
//            s_axis_w_tvalid = 0;
//            s_axis_w_tlast  = 0;
//            #20; // ���
//        end
//    endtask

//    // ���񣺷�������ͼ��
//    task send_image_frame;
//        begin
//            $display("[Time %0t] Starting Image Transmission (%0dx%0d)...", $time, IMG_WIDTH, IMG_HEIGHT);
//            pixel_idx = 0;
            
//            for (r = 0; r < IMG_HEIGHT; r = r + 1) begin
//                for (c = 0; c < IMG_WIDTH; c = c + 1) begin
//                    s_axis_img_tvalid = 1;
//                    // ����ͼ�����ݣ�ÿ��ͨ��ֵ��ͬ
//                    s_axis_img_tdata = 64'h0807060504030201 + pixel_idx; 
                    
//                    if (r == IMG_HEIGHT-1 && c == IMG_WIDTH-1)
//                        s_axis_img_tlast = 1;
//                    else
//                        s_axis_img_tlast = 0;
                    
//                    // �ȴ� Ready
//                    @(posedge clk);
//                    while (s_axis_img_tready == 0) begin
//                        @(posedge clk);
//                    end
                    
//                    pixel_idx = pixel_idx + 1;
//                end
//            end
            
//            s_axis_img_tvalid = 0;
//            s_axis_img_tlast  = 0;
//            $display("[Time %0t] Image Transmission Done.", $time);
//        end
//    endtask

//    // =========================================================================
//    // 6. ����������
//    // =========================================================================
//    reg image_sent_flag;
//    reg compute_done_flag;
    
//    initial begin
//        // --- ��ʼ�� ---
//        rst_n = 0;
//        s_axis_img_tvalid = 0; s_axis_img_tdata = 0; s_axis_img_tlast = 0;
//        s_axis_w_tvalid = 0;   s_axis_w_tdata = 0;   s_axis_w_tlast = 0;
//        m_axis_res_tready = 1; // ʼ��׼���ý��ս��
//        i_load_weights = 0;
//        i_target_layer = 0;
//        i_start_compute = 0;
//        i_l1_weight_base = 0;
//        i_l2_weight_base = 0;
//        received_pixel_cnt = 0;
//        image_sent_flag = 0;
//        compute_done_flag = 0;

//        // --- ��λ ---
//        #100;
//        rst_n = 1;
//        #50;

//        // ---------------------------------------------------------------------
//        // Step 1: ����Ȩ�� (Load Weights)
//        // ---------------------------------------------------------------------
//        // Layer 1 �� 4 �� Core (ID 0~3)
//        // Layer 2 �� 1 �� Core (ID 4)
        
//        // ���� L1 Core 0 (Pattern 0x10)
//        load_weights_for_target(0, 8'h10);
//        // ���� L1 Core 1 (Pattern 0x20)
//        load_weights_for_target(1, 8'h20);
//        // ���� L1 Core 2 (Pattern 0x30)
//        load_weights_for_target(2, 8'h30);
//        // ���� L1 Core 3 (Pattern 0x40)
//        load_weights_for_target(3, 8'h40);
        
//        // ���� L2 Core (ID 4) (Pattern 0x50)
//        load_weights_for_target(4, 8'h50);

//        $display("[Time %0t] All Weights Loaded.", $time);

//        // ---------------------------------------------------------------------
//        // Step 2: ��ʼ���� (Start Compute)
//        // ---------------------------------------------------------------------
//        #100;
//        i_start_compute = 1;
//        i_l1_weight_base = 0; // ʹ�� BRAM ��ַ 0 ��Ȩ��
//        i_l2_weight_base = 0;

//        // ---------------------------------------------------------------------
//        // Step 3: ����ͼ���� (Send Image)
//        // ---------------------------------------------------------------------
//        // ��������
//        send_image_frame();
//        image_sent_flag = 1;
        
//        // �ȴ�һ��ʱ�������
//        #2000;
        
//        $display("\n[Time %0t] Simulation Complete!", $time);
//        $display("Total Output Pixels Received: %d", received_pixel_cnt);
//        if (received_pixel_cnt == IMG_WIDTH * IMG_HEIGHT)
//            $display("TEST PASS: Pixel count matches.");
//        else
//            $display("TEST FAIL: Pixel count mismatch (Expected %d).", IMG_WIDTH * IMG_HEIGHT);
//        $finish;
//    end

//    // =========================================================================
//    // 7. ������
//    // =========================================================================
//    always @(posedge clk) begin
//        if (m_axis_res_tvalid && m_axis_res_tready) begin
//            // ��ӡǰ�����������ڹ۲�
//            if (received_pixel_cnt < 16) begin
//                $display("[Result] Time=%0t Data=%h Last=%b", $time, m_axis_res_tdata, m_axis_res_tlast);
//            end

//            // ���¼��� (���Թ��ƣ�Saver ����߼��� 4 pixels per beat)
//            // ʵ����Ӧ�ÿ� Saver ������߼������������ 4
//            received_pixel_cnt = received_pixel_cnt + 4;
            
//            // �������ź�
//            if (m_axis_res_tlast) begin
//                $display("[Time %0t] Output TLAST detected!", $time);
//            end
//        end
//    end
    
//    // =========================================================================
//    // 8. ��������ź�
//    // =========================================================================
//    always @(posedge clk) begin
//        if (o_compute_done && !compute_done_flag) begin
//            compute_done_flag = 1;
//            $display("[Time %0t] Compute Done signal asserted!", $time);
//        end
//    end

//endmodule
`timescale 1ns / 1ps

module tb_fpga_top_level_new;

    // =========================================================================
    // 1. ��������
    // =========================================================================
    parameter AXIS_DATA_WIDTH = 64;
    parameter NUM_IN_CHANNELS = 8;
    parameter DATA_WIDTH      = 8;
    parameter ACCUM_WIDTH     = 32;
    parameter FILTER_SIZE     = 3;
    
    // ���������16x16 ͼ��
    parameter IMG_WIDTH       = 16;
    parameter IMG_HEIGHT      = 16;
    parameter BRAM_DEPTH      = 512;
    
    // ������ Beat ����256 ���� / 4 ����ÿBeat = 64 Beats
    localparam TOTAL_BEATS    = (IMG_WIDTH * IMG_HEIGHT) / 4; 

    parameter BEATS_PER_WEIGHT_LINE = (NUM_IN_CHANNELS * 2 * FILTER_SIZE * FILTER_SIZE * DATA_WIDTH) / AXIS_DATA_WIDTH;

    // =========================================================================
    // 2. �źŶ���
    // =========================================================================
    reg clk;
    reg rst_n;
    
    // ͼ������
    reg                       s_axis_img_tvalid;
    wire                      s_axis_img_tready;
    reg [AXIS_DATA_WIDTH-1:0] s_axis_img_tdata;
    reg                       s_axis_img_tlast;
    
    // Ȩ������
    reg                       s_axis_w_tvalid;
    wire                      s_axis_w_tready;
    reg [AXIS_DATA_WIDTH-1:0] s_axis_w_tdata;
    reg                       s_axis_w_tlast;
    
    // ������
    wire                      m_axis_res_tvalid;
    reg                       m_axis_res_tready;
    wire [AXIS_DATA_WIDTH-1:0] m_axis_res_tdata;
    wire [AXIS_DATA_WIDTH/8-1:0] m_axis_res_tkeep;
    wire                      m_axis_res_tlast;
    
    // �����ź�
    reg                       i_load_weights;
    reg [3:0]                 i_target_layer;
    reg                       i_start_compute;
    reg [8:0]                 i_l1_weight_base;
    reg [8:0]                 i_l2_weight_base;
    wire                      o_compute_done;
    
    // ͳ����ȶ�
    integer received_pixel_cnt; // ���ؼ���
    integer beat_cnt;           // ���ݰ�����
    integer error_cnt;          // �������
    integer k, r, c, pixel_idx;
    
    // �ƽ�ο����� (64 �� 64-bit ���)
    reg [63:0] golden_data [0:TOTAL_BEATS-1];

    // =========================================================================
    // 3. DUT ʵ����
    // =========================================================================
    fpga_top_level #(
        .AXIS_DATA_WIDTH(AXIS_DATA_WIDTH),
        .NUM_IN_CHANNELS(NUM_IN_CHANNELS),
        .DATA_WIDTH     (DATA_WIDTH),
        .ACCUM_WIDTH    (ACCUM_WIDTH),
        .FILTER_SIZE    (FILTER_SIZE),
        .IMG_WIDTH      (IMG_WIDTH),
        .IMG_HEIGHT     (IMG_HEIGHT),
        .BRAM_DEPTH     (BRAM_DEPTH)
    ) u_dut (
        .clk(clk),
        .rst_n(rst_n),
        .s_axis_img_tvalid(s_axis_img_tvalid),
        .s_axis_img_tready(s_axis_img_tready),
        .s_axis_img_tdata (s_axis_img_tdata),
        .s_axis_img_tlast (s_axis_img_tlast),
        .s_axis_w_tvalid  (s_axis_w_tvalid),
        .s_axis_w_tready  (s_axis_w_tready),
        .s_axis_w_tdata   (s_axis_w_tdata),
        .s_axis_w_tlast   (s_axis_w_tlast),
        .m_axis_res_tvalid(m_axis_res_tvalid),
        .m_axis_res_tready(m_axis_res_tready),
        .m_axis_res_tdata (m_axis_res_tdata),
        .m_axis_res_tkeep (m_axis_res_tkeep),
        .m_axis_res_tlast (m_axis_res_tlast),
        .i_load_weights   (i_load_weights),
        .i_target_layer   (i_target_layer),
        .i_start_compute  (i_start_compute),
        .i_l1_weight_base (i_l1_weight_base),
        .i_l2_weight_base (i_l2_weight_base),
        .o_compute_done   (o_compute_done)
    );

    // =========================================================================
    // 4. ��ʼ���ƽ����� (Golden Reference Initialization)
    // =========================================================================
    initial begin
        // ʹ�� Python �����������ȷֵ
        golden_data[ 0] = 64'h51494f48453f2b27; golden_data[ 1] = 64'h574f564e544c534b;
        golden_data[ 2] = 64'h5e555c535a525950; golden_data[ 3] = 64'h3630564e61575f56;
        golden_data[ 4] = 64'h92848f817e724e47; golden_data[ 5] = 64'h9c8d9a8b97899486;
        golden_data[ 6] = 64'ha696a394a1919e8f; golden_data[ 7] = 64'h5f56988aab9aa998;
        golden_data[ 8] = 64'hc5b2c2afab9b6b60; golden_data[ 9] = 64'hd0bccdbacbb7c8b4;
        golden_data[10] = 64'hdbc6d8c4d6c1d3bf; golden_data[11] = 64'h7d71c8b5e1cbdec9;
        golden_data[12] = 64'hf2daefd8d3bf8477; golden_data[13] = 64'hfde5fae2f7dff4dd;
        golden_data[14] = 64'hffeeffecffe9ffe7; golden_data[15] = 64'h9687f0d9fff3fff1;
        golden_data[16] = 64'hfffffffffbe39d8e; golden_data[17] = 64'hffffffffffffffff;
        golden_data[18] = 64'hffffffffffffffff; golden_data[19] = 64'hae9dfffdffffffff;
        golden_data[20] = 64'hffffffffffffb6a5; golden_data[21] = 64'hffffffffffffffff;
        golden_data[22] = 64'hffffffffffffffff; golden_data[23] = 64'hc7b3ffffffffffff;
        golden_data[24] = 64'hffffffffffffcfbb; golden_data[25] = 64'hffffffffffffffff;
        golden_data[26] = 64'hffffffffffffffff; golden_data[27] = 64'hdfc9ffffffffffff;
        golden_data[28] = 64'hffffffffffffe8d1; golden_data[29] = 64'hffffffffffffffff;
        golden_data[30] = 64'hffffffffffffffff; golden_data[31] = 64'hf7dfffffffffffff;
        golden_data[32] = 64'hffffffffffffffe8; golden_data[33] = 64'hffffffffffffffff;
        golden_data[34] = 64'hffffffffffffffff; golden_data[35] = 64'hfff5ffffffffffff;
        golden_data[36] = 64'hffffffffffffffff; golden_data[37] = 64'hffffffffffffffff;
        golden_data[38] = 64'hffffffffffffffff; golden_data[39] = 64'hffffffffffffffff;
        golden_data[40] = 64'hffffffffffffffff; golden_data[41] = 64'hffffffffffffffff;
        golden_data[42] = 64'hffffffffffffffff; golden_data[43] = 64'hffffffffffffffff;
        golden_data[44] = 64'hffffffffffffffff; golden_data[45] = 64'hffffffffffffffff;
        golden_data[46] = 64'hffffffffffffffff; golden_data[47] = 64'hffffffffffffffff;
        golden_data[48] = 64'hffffffffffffffff; golden_data[49] = 64'hffffffffffffffff;
        golden_data[50] = 64'hffffffffffffffff; golden_data[51] = 64'hffffffffffffffff;
        golden_data[52] = 64'hffffffffffffffff; golden_data[53] = 64'hffffffffffffffff;
        golden_data[54] = 64'hffffffffffffffff; golden_data[55] = 64'hffffffffffffffff;
        golden_data[56] = 64'hffffffffffffffff; golden_data[57] = 64'hffffffffffffffff;
        golden_data[58] = 64'hffffffffffffffff; golden_data[59] = 64'hffffffffffffffff;
        golden_data[60] = 64'hffffffffffffddc7; golden_data[61] = 64'hffffffffffffffff;
        golden_data[62] = 64'hffffffffffffffff; golden_data[63] = 64'hbfacffffffffffff;
    end

    // =========================================================================
    // 5. ʱ������
    // =========================================================================
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    // =========================================================================
    // 6. �������� (Tasks)
    // =========================================================================
    task load_weights_for_target;
        input [3:0] target_id;
        input [7:0] start_val;
        reg [7:0] k_val;
        begin
            $display("[Time %0t] Loading Weights for Target ID: %d", $time, target_id);
            @(posedge clk);
            i_target_layer = target_id;
            i_load_weights = 1;
            @(posedge clk);
            i_load_weights = 0;
            
            for (k = 0; k < BEATS_PER_WEIGHT_LINE; k = k + 1) begin
                s_axis_w_tvalid = 1;
                k_val = start_val + k;
                s_axis_w_tdata  = {8{k_val}};
                s_axis_w_tlast  = (k == BEATS_PER_WEIGHT_LINE - 1);
                @(posedge clk);
            end
            s_axis_w_tvalid = 0;
            s_axis_w_tlast  = 0;
            #20;
        end
    endtask

    task send_image_frame;
        begin
            $display("[Time %0t] Starting Image Transmission (%0dx%0d)...", $time, IMG_WIDTH, IMG_HEIGHT);
            pixel_idx = 0;
            for (r = 0; r < IMG_HEIGHT; r = r + 1) begin
                for (c = 0; c < IMG_WIDTH; c = c + 1) begin
                    s_axis_img_tvalid = 1;
                    s_axis_img_tdata = 64'h0807060504030201 + pixel_idx;
                    s_axis_img_tlast = (r == IMG_HEIGHT-1 && c == IMG_WIDTH-1);
                    @(posedge clk);
                    while (s_axis_img_tready == 0) @(posedge clk);
                    pixel_idx = pixel_idx + 1;
                end
            end
            s_axis_img_tvalid = 0;
            s_axis_img_tlast  = 0;
            $display("[Time %0t] Image Transmission Done.", $time);
        end
    endtask

    // =========================================================================
    // 7. ������
    // =========================================================================
    reg [31:0] watchdog;
    
    initial begin
        // --- ��ʼ�� ---
        rst_n = 0;
        s_axis_img_tvalid = 0; s_axis_img_tdata = 0; s_axis_img_tlast = 0;
        s_axis_w_tvalid = 0;   s_axis_w_tdata = 0;   s_axis_w_tlast = 0;
        m_axis_res_tready = 1; 
        i_load_weights = 0; i_target_layer = 0; i_start_compute = 0;
        i_l1_weight_base = 0; i_l2_weight_base = 0;
        received_pixel_cnt = 0;
        beat_cnt = 0;
        error_cnt = 0;
        
        // --- ��λ ---
        #100; rst_n = 1; #50;

        // Step 1: ����Ȩ��
        load_weights_for_target(0, 8'h10);
        load_weights_for_target(1, 8'h20);
        load_weights_for_target(2, 8'h30);
        load_weights_for_target(3, 8'h40);
        load_weights_for_target(4, 8'h50);

        // Step 2: ��������
        #100;
        i_start_compute = 1;

        // Step 3: ����ͼ��
        send_image_frame();

        // Step 4: �ȴ����
        $display("[Time %0t] Waiting for results...", $time);
        watchdog = 0;
        while (received_pixel_cnt < IMG_WIDTH * IMG_HEIGHT && watchdog < 10000) begin
            @(posedge clk);
            watchdog = watchdog + 1;
        end
        
        #100;
        $display("\n=================================================");
        $display("          SIMULATION REPORT");
        $display("=================================================");
        $display("Total Beats Received: %d / %d", beat_cnt, TOTAL_BEATS);
        $display("Total Pixels: %d / %d", received_pixel_cnt, IMG_WIDTH*IMG_HEIGHT);
        
        if (error_cnt == 0 && beat_cnt == TOTAL_BEATS) begin
            $display("\n[SUCCESS] ALL DATA MATCHED GOLDEN REFERENCE!");
        end else begin
            $display("\n[FAILURE] Found %d Mismatches.", error_cnt);
            if (beat_cnt != TOTAL_BEATS)
                $display("[FAILURE] Data count mismatch (Expected %d beats).", TOTAL_BEATS);
        end
        $display("=================================================");
        $stop;
    end

    // =========================================================================
    // 8. ��������ȶ� (Monitor & Checker)
    // =========================================================================
    always @(posedge clk) begin
        if (m_axis_res_tvalid && m_axis_res_tready) begin
            // ��ӡ���ȶ�
            if (beat_cnt < TOTAL_BEATS) begin
                if (m_axis_res_tdata === golden_data[beat_cnt]) begin
                    $display("[CHECK PASS] Beat %2d: Data=%h (Matched)", beat_cnt, m_axis_res_tdata);
                end else begin
                    $display("[CHECK FAIL] Beat %2d: Data=%h | Exp=%h !!!", beat_cnt, m_axis_res_tdata, golden_data[beat_cnt]);
                    error_cnt = error_cnt + 1;
                end
            end else begin
                $display("[WARNING] Received extra beat: %h", m_axis_res_tdata);
            end

            // ���¼�����
            beat_cnt = beat_cnt + 1;
            received_pixel_cnt = received_pixel_cnt + 4; // ÿ�� Beat 4 �����أ�ÿ������ 2 �����ͨ��? 
            // ����������֮ǰ�ķ�����һ��Beat�� 4 ������ (64bit / 16bit_per_pixel)
            // �����������ؼ���Ӧ���� +4�������� +8��
            // �������� Saver ������ÿ��ʱ�ӳ� 8 ��ͨ�����Ǿ��� +8��
            // �����Ǳ��ֺ�֮ǰ����һ�µ� +4 (4 pixels * 2 channels * 8 bits = 64 bits)
            
            if (m_axis_res_tlast) begin
                $display("[Time %0t] TLAST detected!", $time);
            end
        end
    end

endmodule