`timescale 1ns / 1ps

module dynamic_line_buffer #(
    parameter DATA_WIDTH = 8,
    parameter MAX_DEPTH  = 2048  // ֧�ֵ����ͼ����
)(
    input                       clk,
    input                       rst_n,
    
    input                       i_valid,       // дʹ��
    input  [15:0]               i_width,       // ���ؼ�����ǰͼ����
    input  [DATA_WIDTH-1:0]     i_data,        // ��������
    output [DATA_WIDTH-1:0]     o_data         // ������� (�ӳ���һ�е�����)
);

    // --- ָ�붨�� ---
    // ʹ�ñ� log2(MAX_DEPTH) ��һλ��λ�����㴦��ָ����ƺͼ���
    reg [$clog2(MAX_DEPTH):0]   wr_ptr;
    wire [$clog2(MAX_DEPTH):0]  rd_ptr_calc;
    
    // ʵ�� RAM ��ַ
    wire [$clog2(MAX_DEPTH)-1:0] wr_addr;
    wire [$clog2(MAX_DEPTH)-1:0] rd_addr;

    // --- 1. дָ���߼� (�򵥵Ļ��μ���) ---
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            wr_ptr <= 0;
        end else if (i_valid) begin
            if (wr_ptr == MAX_DEPTH - 1)
                wr_ptr <= 0;
            else
                wr_ptr <= wr_ptr + 1;
        end
    end

    // --- 2. ����ַ���� (�����������ӳٲ���) ---
    // ԭ��BRAM ��ȡ������Ҫ 1 ��ʱ�����ڡ�
    // ������������������ o_data �뵱ǰ���� i_data ���߼���������� i_width �����ڣ�
    // ���Ǳ���"��ǰ"һ��λ�ö�ȡ������ BRAM �Ķ��ӳ١�
    // Read_Ptr = Write_Ptr - (Width - 1)
    
    wire [$clog2(MAX_DEPTH):0] latency_offset;
    assign latency_offset = i_width - 1; 

    // �����λ������ļ�������
    assign rd_ptr_calc = (wr_ptr >= latency_offset) ? 
                         (wr_ptr - latency_offset) : 
                         (wr_ptr + MAX_DEPTH - latency_offset);
    
    assign wr_addr = wr_ptr[$clog2(MAX_DEPTH)-1:0];
    assign rd_addr = rd_ptr_calc[$clog2(MAX_DEPTH)-1:0];

    // --- 3. �ƶ�˫�˿� RAM (Inferred BRAM) ---
    reg [DATA_WIDTH-1:0] ram [0:MAX_DEPTH-1];
    reg [DATA_WIDTH-1:0] ram_out;

    always @(posedge clk) begin
        if (i_valid) begin
            ram[wr_addr] <= i_data;
        end
    end

    always @(posedge clk) begin
        // ֻҪʱ�����ܣ��ͳ�����ȡ��һ�е�����
        // �����Ҫ���ϸ�Ĺ��Ŀ��ƣ����Խ� i_valid ��Ϊ��ʹ��
        ram_out <= ram[rd_addr]; 
    end

    assign o_data = ram_out;

endmodule