`timescale 1ns / 1ps

module feature_map_saver_axis #(
    parameter AXIS_DATA_WIDTH = 64,      // DMA �ӿ�λ��
    parameter INPUT_WIDTH     = 35,      // ��������λ�� (���� 32λ�ۼ� + log2(8ͨ��) �� 35)
    parameter OUTPUT_WIDTH    = 8,       // �����DDR��λ�� (uint8)
    parameter QUANT_SHIFT     = 10       // ��������λ�� (�൱�ڳ��� 2^10)
)(
    input                               clk,
    input                               rst_n,

    // =========================================================================
    // 1. ���� Conv Core ������ӿ�
    // =========================================================================
    input                               i_valid,
    input        signed [INPUT_WIDTH-1:0] i_data_A, // Kernel A �Ľ�� (ͨ�� N)
    input        signed [INPUT_WIDTH-1:0] i_data_B, // Kernel B �Ľ�� (ͨ�� N+1)
    
    // =========================================================================
    // 2. ͼ����� (�������� TLAST)
    // =========================================================================
    // ͼ���������� = Height * Width (�ռ�������������ͨ��)
    // ģ����Զ����ݴ���߼������ʱ���� TLAST
    input        [31:0]                 i_total_pixels, 
    
    // =========================================================================
    // 3. AXI-Stream Master ��� (���� DMA S2MM)
    // =========================================================================
    output reg                          m_axis_tvalid,
    input                               m_axis_tready,
    output reg   [AXIS_DATA_WIDTH-1:0]  m_axis_tdata,
    output reg   [AXIS_DATA_WIDTH/8-1:0]m_axis_tkeep,
    output reg                          m_axis_tlast
);

    // =========================================================================
    // Stage 1: ���� (ReLU + Quantization + Clamp)
    // =========================================================================
    reg [OUTPUT_WIDTH-1:0] post_data_A;
    reg [OUTPUT_WIDTH-1:0] post_data_B;
    reg                    post_valid;

    // ����������
    function [OUTPUT_WIDTH-1:0] process_pixel;
        input signed [INPUT_WIDTH-1:0] raw_in;
        reg signed [INPUT_WIDTH-1:0] shifted;
        begin
            // 1. ReLU: ������0
            if (raw_in < 0) begin
                process_pixel = 0;
            end else begin
                // 2. Scaling: �������� (�൱�ڳ��� 2^QUANT_SHIFT)
                shifted = raw_in >>> QUANT_SHIFT;
                
                // 3. Clamping: ���ͽضϵ� 8-bit (0~255)
                // ����Ƿ񳬹����ֵ (2^8 - 1 = 255)
                if (shifted > { {(INPUT_WIDTH-OUTPUT_WIDTH){1'b0}}, {(OUTPUT_WIDTH){1'b1}} }) 
                    process_pixel = {(OUTPUT_WIDTH){1'b1}}; // 255
                else
                    process_pixel = shifted[OUTPUT_WIDTH-1:0];
            end
        end
    endfunction

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            post_valid <= 0;
            post_data_A <= 0;
            post_data_B <= 0;
        end else begin
            post_valid <= i_valid;
            if (i_valid) begin
                post_data_A <= process_pixel(i_data_A);
                post_data_B <= process_pixel(i_data_B);
            end
        end
    end

    // =========================================================================
    // Stage 2: ���ݴ�� (Packing)
    // =========================================================================
    // Ŀ�꣺��ÿ������� 2 �� 8-bit ����ƴ�ճ� 64-bit ��������
    // ��Ҫ���� 4 ����Ч����������� 64-bit (2 bytes * 4 = 8 bytes)
    
    reg [AXIS_DATA_WIDTH-1:0] pack_buffer; // ��λ�Ĵ���/����
    reg [1:0]                 pack_cnt;    // ������ 0..3
    
    // TLAST ���ؼ�����
    reg [31:0]                pixel_counter;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            m_axis_tvalid <= 0;
            m_axis_tdata  <= 0;
            m_axis_tkeep  <= 8'hFF;
            m_axis_tlast  <= 0;
            pack_cnt      <= 0;
            pack_buffer   <= 0;
            pixel_counter <= 0;
        end else begin
            // �����߼�������ӻ�Ready�������Valid��׼����һ�δ���
            if (m_axis_tready && m_axis_tvalid) begin
                m_axis_tvalid <= 0;
                m_axis_tlast  <= 0;
            end

            if (post_valid) begin
                // ���� Buffer: ���� Little-Endian (�͵�ַ�ŵ�λ)
                // ÿ������ 16 bits (Data B @ High, Data A @ Low)
                // pack_cnt=0: [15:0], pack_cnt=1: [31:16], ...
                pack_buffer[pack_cnt*16 +: 16] <= {post_data_B, post_data_A};
                
                // �������ؼ��� (ÿ�� valid ʱ�Ӵ��� 1 ���ռ�λ��)
                if (pixel_counter < i_total_pixels - 1)
                    pixel_counter <= pixel_counter + 1;
                else
                    pixel_counter <= 0;

                // -------------------------------------------------------------
                // ���������ж�
                // -------------------------------------------------------------
                // 1. Buffer ������ (pack_cnt == 3)
                // 2. ���� �Ѿ������һ�������� (��Ҫǿ�Ʒ���ʣ��Ĳ�������)
                if (pack_cnt == 3 || pixel_counter == i_total_pixels - 1) begin
                    
                    m_axis_tvalid <= 1;
                    
                    // ����ǰ����ƴ�ӵ� buffer ��λ�����
                    // ע�⣺pack_buffer �д洢����ǰ 0~2 �ε����ݣ���ǰ�� 3 �ε�����ֱ��������
                    // �����λ���߼�ȷ������˳����ȷ��D3_D2_D1_D0 (D0�ڵ�λ)
                    // ��������һ�δ����� pack_cnt < 3����Ҫ���⴦�����ݶ���
                    
                    case (pack_cnt)
                        0: m_axis_tdata <= { {(64-16){1'b0}}, post_data_B, post_data_A };
                        1: m_axis_tdata <= { {(64-32){1'b0}}, post_data_B, post_data_A, pack_buffer[15:0] };
                        2: m_axis_tdata <= { {(64-48){1'b0}}, post_data_B, post_data_A, pack_buffer[31:0] };
                        3: m_axis_tdata <= { post_data_B, post_data_A, pack_buffer[47:0] };
                    endcase
                    
                    // ���� TLAST �� TKEEP
                    if (pixel_counter == i_total_pixels - 1) begin
                        m_axis_tlast <= 1;
                        // ������Ч�ֽ� (Strobe)
                        // pack_cnt=0 -> 2 bytes, =1 -> 4 bytes, =2 -> 6 bytes, =3 -> 8 bytes
                        case(pack_cnt)
                            0: m_axis_tkeep <= 8'b0000_0011;
                            1: m_axis_tkeep <= 8'b0000_1111;
                            2: m_axis_tkeep <= 8'b0011_1111;
                            3: m_axis_tkeep <= 8'b1111_1111;
                        endcase
                        pack_cnt <= 0; // ֡������λ
                    end else begin
                        m_axis_tlast <= 0;
                        m_axis_tkeep <= 8'hFF; // �м�����ȫ��Ч
                        pack_cnt <= 0;         // ������λ
                    end
                end else begin
                    // ��û���Ҳ������һ����������
                    pack_cnt <= pack_cnt + 1;
                end
            end
        end
    end

endmodule