`timescale 1ns / 1ps

module tb_fpga_top_level;

    // =========================================================================
    // 1. ��������
    // =========================================================================
    parameter AXIS_DATA_WIDTH = 64;
    parameter NUM_IN_CHANNELS = 8;
    parameter DATA_WIDTH      = 8;
    parameter ACCUM_WIDTH     = 32;
    parameter FILTER_SIZE     = 3;
    
    // Ϊ�˷����ٶȣ����ǽ�ͼ��ߴ���Сһ��
    parameter IMG_WIDTH       = 16; 
    parameter IMG_HEIGHT      = 16;
    parameter BRAM_DEPTH      = 512;

    // Ȩ�ؼ�����ؼ���
    // Layer 1: 4 Cores, ÿ�� Core ���� 2 �����ͨ��
    // ÿ�� Core ��Ҫ 144 ��Ȩ�� (8 In * 2 Out * 9) = 1152 bits
    // 1152 bits / 64 bits (AXI) = 18 Beats
    localparam BEATS_PER_WEIGHT_LINE = (NUM_IN_CHANNELS * 2 * FILTER_SIZE * FILTER_SIZE * DATA_WIDTH) / AXIS_DATA_WIDTH;

    // =========================================================================
    // 2. �źŶ���
    // =========================================================================
    reg clk;
    reg rst_n;

    // ͼ������
    reg                       s_axis_img_tvalid;
    wire                      s_axis_img_tready;
    reg [AXIS_DATA_WIDTH-1:0] s_axis_img_tdata;
    reg                       s_axis_img_tlast;

    // Ȩ������
    reg                       s_axis_w_tvalid;
    wire                      s_axis_w_tready;
    reg [AXIS_DATA_WIDTH-1:0] s_axis_w_tdata;
    reg                       s_axis_w_tlast;

    // ������
    wire                      m_axis_res_tvalid;
    reg                       m_axis_res_tready;
    wire [AXIS_DATA_WIDTH-1:0] m_axis_res_tdata;
    wire [AXIS_DATA_WIDTH/8-1:0] m_axis_res_tkeep;
    wire                      m_axis_res_tlast;

    // �����ź�
    reg                       i_load_weights;
    reg [3:0]                 i_target_layer;
    reg                       i_start_compute;
    reg [8:0]                 i_l1_weight_base;
    reg [8:0]                 i_l2_weight_base;
    wire                      o_compute_done;

    assign s_axis_w_tready = 1'b1;
    // ͳ�ƽ��յ���������
    integer received_pixel_cnt;

    // =========================================================================
    // 3. DUT ʵ����
    // =========================================================================
    fpga_top_level #(
        .AXIS_DATA_WIDTH(AXIS_DATA_WIDTH),
        .NUM_IN_CHANNELS(NUM_IN_CHANNELS),
        .DATA_WIDTH     (DATA_WIDTH),
        .ACCUM_WIDTH    (ACCUM_WIDTH),
        .FILTER_SIZE    (FILTER_SIZE),
        .IMG_WIDTH      (IMG_WIDTH),
        .IMG_HEIGHT     (IMG_HEIGHT),
        .BRAM_DEPTH     (BRAM_DEPTH)
    ) u_dut (
        .clk(clk),
        .rst_n(rst_n),
        
        .s_axis_img_tvalid(s_axis_img_tvalid),
        .s_axis_img_tready(s_axis_img_tready),
        .s_axis_img_tdata (s_axis_img_tdata),
        .s_axis_img_tlast (s_axis_img_tlast),
        
        .s_axis_w_tvalid  (s_axis_w_tvalid),
        .s_axis_w_tready  (s_axis_w_tready),
        .s_axis_w_tdata   (s_axis_w_tdata),
        .s_axis_w_tlast   (s_axis_w_tlast),
        
        .m_axis_res_tvalid(m_axis_res_tvalid),
        .m_axis_res_tready(m_axis_res_tready),
        .m_axis_res_tdata (m_axis_res_tdata),
        .m_axis_res_tkeep (m_axis_res_tkeep),
        .m_axis_res_tlast (m_axis_res_tlast),
        
        .i_load_weights   (i_load_weights),
        .i_target_layer   (i_target_layer),
        .i_start_compute  (i_start_compute),
        .i_l1_weight_base (i_l1_weight_base),
        .i_l2_weight_base (i_l2_weight_base),
        .o_compute_done   (o_compute_done)
    );

    // =========================================================================
    // 4. ʱ������ (100MHz)
    // =========================================================================
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    // =========================================================================
    // 5. ������ (Helper Tasks)
    // =========================================================================
    
    // ���񣺼���һ��Ȩ�ص�ָ���� Target Layer
    task load_weights_for_target(input [3:0] target_id, input [7:0] start_val);
        integer k;
        begin
            $display("[Time %0t] Loading Weights for Target ID: %d", $time, target_id);
            
            // 1. ���ÿ����ź�
            @(posedge clk);
            i_target_layer = target_id;
            i_load_weights = 1; // ������λ����
            @(posedge clk);
            i_load_weights = 0; // �������壬��ʼ����
            
            // 2. ���� AXI Stream ����
            // ����ÿ�� Core ֻ��Ҫ 1 ��Ȩ�� (Addr 0)����Ҫ���� BEATS_PER_WEIGHT_LINE ��
            for (k = 0; k < BEATS_PER_WEIGHT_LINE; k = k + 1) begin
                s_axis_w_tvalid = 1;
                // ����������ݣ��򵥵ĵ��������������
                s_axis_w_tdata  = {8{start_val + k[7:0]}}; 
                
                if (k == BEATS_PER_WEIGHT_LINE - 1) 
                    s_axis_w_tlast = 1;
                else 
                    s_axis_w_tlast = 0;
                
                @(posedge clk);
            end
            
            s_axis_w_tvalid = 0;
            s_axis_w_tlast  = 0;
            #20; // ���
        end
    endtask

    // ���񣺷�������ͼ��
// ���񣺷�������ͼ��
    task send_image_frame();
        integer r, c;
        integer pixel_idx;
        begin
            $display("[Time %0t] Starting Image Transmission (%0dx%0d)...", $time, IMG_WIDTH, IMG_HEIGHT);
            pixel_idx = 0;
            
            for (r = 0; r < IMG_HEIGHT; r = r + 1) begin
                for (c = 0; c < IMG_WIDTH; c = c + 1) begin
                    s_axis_img_tvalid = 1;
                    // ����ͼ�����ݣ�ÿ��ͨ��ֵ��ͬ
                    s_axis_img_tdata = 64'h0807060504030201 + pixel_idx; 
                    
                    if (r == IMG_HEIGHT-1 && c == IMG_WIDTH-1)
                        s_axis_img_tlast = 1;
                    else
                        s_axis_img_tlast = 0;
                    
                    // --- �������ֿ�ʼ ---
                    // �ȴ� Ready (��׼ Verilog д��)
                    @(posedge clk);
                    while (!s_axis_img_tready) begin
                        @(posedge clk);
                    end
                    // --- �������ֽ��� ---
                    
                    pixel_idx = pixel_idx + 1;
                end
            end
            
            s_axis_img_tvalid = 0;
            s_axis_img_tlast  = 0;
            $display("[Time %0t] Image Transmission Done.", $time);
        end
    endtask

    // =========================================================================
    // 6. ����������
    // =========================================================================
    initial begin
        // --- ��ʼ�� ---
        rst_n = 0;
        s_axis_img_tvalid = 0; s_axis_img_tdata = 0; s_axis_img_tlast = 0;
        s_axis_w_tvalid = 0;   s_axis_w_tdata = 0;   s_axis_w_tlast = 0;
        m_axis_res_tready = 1; // ʼ��׼���ý��ս��
        i_load_weights = 0;
        i_target_layer = 0;
        i_start_compute = 0;
        i_l1_weight_base = 0;
        i_l2_weight_base = 0;
        received_pixel_cnt = 0;

        // --- ��λ ---
        #100;
        rst_n = 1;
        #50;

        // ---------------------------------------------------------------------
        // Step 1: ����Ȩ�� (Load Weights)
        // ---------------------------------------------------------------------
        // Layer 1 �� 4 �� Core (ID 0~3)
        // Layer 2 �� 1 �� Core (ID 4)
        
        // ���� L1 Core 0 (Pattern 0x10)
        load_weights_for_target(0, 8'h10);
        // ���� L1 Core 1 (Pattern 0x20)
        load_weights_for_target(1, 8'h20);
        // ���� L1 Core 2 (Pattern 0x30)
        load_weights_for_target(2, 8'h30);
        // ���� L1 Core 3 (Pattern 0x40)
        load_weights_for_target(3, 8'h40);
        
        // ���� L2 Core (ID 4) (Pattern 0x50)
        load_weights_for_target(4, 8'h50);

        $display("[Time %0t] All Weights Loaded.", $time);

        // ---------------------------------------------------------------------
        // Step 2: ��ʼ���� (Start Compute)
        // ---------------------------------------------------------------------
        #100;
        i_start_compute = 1;
        i_l1_weight_base = 0; // ʹ�� BRAM ��ַ 0 ��Ȩ��
        i_l2_weight_base = 0;

        // ---------------------------------------------------------------------
        // Step 3: ����ͼ���� (Send Image)
        // ---------------------------------------------------------------------
        fork
            // �߳� 1: ��������
            send_image_frame();
            
            // �߳� 2: �������ź�
            begin
                wait(o_compute_done);
                $display("\n[Time %0t] Compute Done Interrupt Received!", $time);
                #100;
                $display("Total Output Pixels Received: %d", received_pixel_cnt);
                if (received_pixel_cnt == IMG_WIDTH * IMG_HEIGHT)
                    $display("TEST PASS: Pixel count matches.");
                else
                    $display("TEST FAIL: Pixel count mismatch (Expected %d).", IMG_WIDTH * IMG_HEIGHT);
                $finish;
            end
        join
    end

    // =========================================================================
    // 7. ������
    // =========================================================================
    always @(posedge clk) begin
        if (m_axis_res_tvalid && m_axis_res_tready) begin
            // ����� pack_cnt �߼�ȡ���� Saver ģ�飬ÿ 4 �����س�һ�� 64bit
            // �� Saver �ڲ��� pixel_counter �ǰ����ؼ�����
            // ����������Ǽ��� tvalid ÿ����һ�Σ������� 4 ������ (�������һ�ο�����)
            
            // ��ӡǰ�����������ڹ۲�
            if (received_pixel_cnt < 16) begin
                $display("[Result] Time=%0t Data=%h Last=%b", $time, m_axis_res_tdata, m_axis_res_tlast);
            end

            // ���¼��� (���Թ��ƣ�Saver ����߼��� 4 pixels per beat)
            // ʵ����Ӧ�ÿ� Saver ������߼������������ 4
            received_pixel_cnt = received_pixel_cnt + 4;
        end
    end

endmodule