`timescale 1ns / 1ps

module line_buffer_with_padding #(
    parameter NUM_CHANNELS = 8,
    parameter DATA_WIDTH   = 8,
    parameter IMG_WIDTH    = 256,
    parameter IMG_HEIGHT   = 256,
    parameter FILTER_SIZE  = 3
)(
    input                                   clk,
    input                                   rst_n,
    input                                   i_valid,
    input [NUM_CHANNELS*DATA_WIDTH-1:0]     i_data_parallel,
    output reg                              o_valid,
    output [NUM_CHANNELS*FILTER_SIZE*FILTER_SIZE*DATA_WIDTH-1:0] o_windows_packed
);

    localparam TOTAL_DATA_WIDTH = NUM_CHANNELS * DATA_WIDTH;

    // =========================================================================
    // 1. Line Buffers & ·��ƽ�� (Path Balancing)
    // =========================================================================
    // Ŀ�꣺��� BRAM �ۻ��ӳٵ��µĽ��ݴ�λ
    // �ӳٷ�����
    // LB Output Latency = Width + 1 (1 cycle BRAM read)
    // Row 0 (Input): Latency 0
    // Row 1 (LB0)  : Latency W + 1
    // Row 2 (LB1)  : Latency 2W + 2
    
    // ԭʼ���
    wire [TOTAL_DATA_WIDTH-1:0] lb0_out; // ԭʼ LB0 ���
    wire [TOTAL_DATA_WIDTH-1:0] lb1_out; // ԭʼ LB1 ��� (Top Row, ����)

    // ������������
    reg  [TOTAL_DATA_WIDTH-1:0] row_0_aligned; // Bot Row (���ӳ� 2 cycles)
    reg  [TOTAL_DATA_WIDTH-1:0] row_1_aligned; // Mid Row (���ӳ� 1 cycle)
    wire [TOTAL_DATA_WIDTH-1:0] row_2_aligned; // Top Row (��׼����������ӳ�)

    // �����Ĵ������ڴ���
    reg [TOTAL_DATA_WIDTH-1:0] row_0_d1; 

    // --- Line Buffer ʵ���� ---
    dynamic_line_buffer #(.DATA_WIDTH(TOTAL_DATA_WIDTH), .MAX_DEPTH(IMG_WIDTH)) u_lb0 (
        .clk(clk), .i_valid(i_valid), .i_width(IMG_WIDTH[15:0]), 
        .i_data(i_data_parallel), .o_data(lb0_out)
    );

    dynamic_line_buffer #(.DATA_WIDTH(TOTAL_DATA_WIDTH), .MAX_DEPTH(IMG_WIDTH)) u_lb1 (
        .clk(clk), .i_valid(i_valid), .i_width(IMG_WIDTH[15:0]), 
        .i_data(lb0_out),         .o_data(lb1_out)
    );

    // --- �ؼ���Ӳ�����Ķ��� ---
    always @(posedge clk) begin
        if (i_valid) begin
            // Row 0 (Bot): Input -> Delay 1 -> Delay 2
            row_0_d1      <= i_data_parallel;
            row_0_aligned <= row_0_d1;      // �ӳ� 2 �ģ����� Top
            
            // Row 1 (Mid): LB0_Out -> Delay 1
            row_1_aligned <= lb0_out;       // �ӳ� 1 �ģ����� Top
        end
    end
    
    // Row 2 (Top): ֱ��ʹ�ã���Ϊ���������� (�ӳ� 2 ������ 2��BRAM)
    assign row_2_aligned = lb1_out;

    // =========================================================================
    // 2. ��λ�Ĵ��� (Shift Register)
    // =========================================================================
    reg [DATA_WIDTH-1:0] window_raw [NUM_CHANNELS-1:0][FILTER_SIZE-1:0][FILTER_SIZE-1:0];
    integer c;
    
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            // reset
        end else if (i_valid) begin
            for (c = 0; c < NUM_CHANNELS; c = c + 1) begin
                // Row 0 (Top) <--- row_2_aligned (��ɵ�����)
                window_raw[c][0][0] <= window_raw[c][0][1];
                window_raw[c][0][1] <= window_raw[c][0][2];
                window_raw[c][0][2] <= row_2_aligned[c*DATA_WIDTH +: DATA_WIDTH];
                
                // Row 1 (Mid) <--- row_1_aligned
                window_raw[c][1][0] <= window_raw[c][1][1];
                window_raw[c][1][1] <= window_raw[c][1][2];
                window_raw[c][1][2] <= row_1_aligned[c*DATA_WIDTH +: DATA_WIDTH];

                // Row 2 (Bot) <--- row_0_aligned (�������ݣ����ӳٶ���)
                window_raw[c][2][0] <= window_raw[c][2][1];
                window_raw[c][2][1] <= window_raw[c][2][2];
                window_raw[c][2][2] <= row_0_aligned[c*DATA_WIDTH +: DATA_WIDTH];
            end
        end
    end

    // =========================================================================
    // 3. ������ Valid ����
    // =========================================================================
    reg [15:0] col_ptr;
    reg [15:0] row_ptr;
    
    // �������������ͺ��� 2 ������ (���뵽��������·��)��
    // ��Ч�����ĵ����Ҳ��Ҫ��Ӧƥ�䡣
    // ����Ϊ col_ptr Ҳ������ i_valid ���µģ�������ͬ���ƽ��ġ�
    // ����ֻ��Ҫ��֤ padding �߼����õ���"��ǰ�� shift register ����"�����꼴�ɡ�
    
    wire signed [16:0] center_x = col_ptr - 1;
    wire signed [16:0] center_y = row_ptr - 1;
    reg pad_top, pad_bottom, pad_left, pad_right;
    reg center_valid;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            col_ptr <= 0; row_ptr <= 0;
            pad_top <= 0; pad_bottom <= 0; pad_left <= 0; pad_right <= 0;
            center_valid <= 0;
        end else if (i_valid) begin
            // �������
            if (col_ptr == IMG_WIDTH - 1) begin
                col_ptr <= 0;
                if (row_ptr == IMG_HEIGHT - 1) row_ptr <= 0;
                else row_ptr <= row_ptr + 1;
            end else begin
                col_ptr <= col_ptr + 1;
            end

            // Padding ��־
            pad_top    <= (center_y == 0);
            pad_bottom <= (center_y == IMG_HEIGHT - 1);
            pad_left   <= (center_x == 0);
            pad_right  <= (center_x == IMG_WIDTH - 1);

            // Valid �ж�
            // �������ӳٶ����������Ҫ�ȴ� LineBuffer ������
            // ��Ȼ�ǵȴ��� 1 �� (row_ptr=1) ��ʼ����ʱ�����ܲ�����Ч����
            if (row_ptr == 0)
                center_valid <= 0;
            else
                center_valid <= 1;

        end else begin
            // ����Ҫ��������Чʱ���������� valid����ֹ��ѭ��
            center_valid <= 0;
        end
    end
    
    // ��� Valid ��һ�ģ�ƥ�� Shift Register ���������
    always @(posedge clk) o_valid <= center_valid;

    // =========================================================================
    // 4. ������
    // =========================================================================
    genvar gc, gr, gk;
    generate
        for (gc = 0; gc < NUM_CHANNELS; gc = gc + 1) begin : loop_ch
            for (gr = 0; gr < FILTER_SIZE; gr = gr + 1) begin : loop_row
                for (gk = 0; gk < FILTER_SIZE; gk = gk + 1) begin : loop_col
                    wire is_masked = (pad_top && (gr == 0)) || (pad_bottom && (gr == 2)) ||
                                     (pad_left && (gk == 0)) || (pad_right  && (gk == 2));
                    wire [DATA_WIDTH-1:0] raw = window_raw[gc][gr][gk];
                    assign o_windows_packed[(gc*9 + gr*3 + gk)*DATA_WIDTH +: DATA_WIDTH] = 
                           is_masked ? {DATA_WIDTH{1'b0}} : raw;
                end
            end
        end
    endgenerate

endmodule