module simple_dual_port_ram_dynamic #(parameter WIDTH=8, DEPTH=512)(
    input clk, input we, 
    input [$clog2(DEPTH)-1:0] wr_addr, rd_addr,
    input [WIDTH-1:0] din, output reg [WIDTH-1:0] dout
);
    (* ram_style = "block" *) reg [WIDTH-1:0] ram [0:DEPTH-1];
    
    // ��ʼ�� RAM �Ա�����治��̬ (��ѡ)
    integer i;
    initial begin
        for(i=0; i<DEPTH; i=i+1) ram[i] = 0;
    end

    always @(posedge clk) begin
        if (we) ram[wr_addr] <= din;
        dout <= ram[rd_addr]; // ���ӳ� 1 ��
    end
endmodule
