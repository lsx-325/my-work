`timescale 1ns / 1ps

module axis_ping_pong_buffer #(
    parameter DATA_WIDTH = 64,
    parameter ADDR_WIDTH = 6,   // 2^6 = 64 depth
    parameter MAX_DEPTH  = 64
)(
    input  wire                   clk,
    input  wire                   rst_n,

    // ========================================
    // AXI-Stream Slave (Input / Upstream)
    // ========================================
    input  wire [DATA_WIDTH-1:0]  s_axis_tdata,
    input  wire                   s_axis_tvalid,
    input  wire                   s_axis_tlast,
    output wire                   s_axis_tready,

    // ========================================
    // AXI-Stream Master (Output / Downstream)
    // ========================================
    output reg  [DATA_WIDTH-1:0]  m_axis_tdata,
    output reg                    m_axis_tvalid,
    output reg                    m_axis_tlast,
    input  wire                   m_axis_tready
);

    // =========================================================================
    // 1. �ڴ涨�� (Distributed RAM �� Block RAM ������)
    // =========================================================================
    reg [DATA_WIDTH-1:0] ram_buf0 [0:MAX_DEPTH-1];
    reg [DATA_WIDTH-1:0] ram_buf1 [0:MAX_DEPTH-1];

    // ���ȱ��붨��Ϊ ADDR_WIDTH + 1 λ�����ܹ��洢��ֵ "64"
    reg [ADDR_WIDTH:0]   len_buf0, len_buf1; 

    // Buffer ״̬: 0 = ��/����д, 1 = ��/����ȡ
    reg [1:0] buf_full; 

    // =========================================================================
    // 2. д���߼� (Write Control)
    // =========================================================================
    reg [ADDR_WIDTH:0] wr_ptr;      
    reg                wr_sel;      // ��ǰ����д�� buffer ���� (0/1)
    
    // ֻ�е���ǰѡ�е� buffer ����ʱ������Ϊ�������ṩ Ready
    assign s_axis_tready = !buf_full[wr_sel];

    wire wr_handshake = s_axis_tvalid && s_axis_tready;
    wire wr_finish    = wr_handshake && (s_axis_tlast || (wr_ptr == MAX_DEPTH-1));

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            wr_ptr   <= 0;
            wr_sel   <= 0;
            buf_full <= 2'b00;
            len_buf0 <= 0;
            len_buf1 <= 0;
        end else begin
            // --- ״̬��� ---
            // ���ն�ȡ��������źţ���� Full ��־
            if (rd_buf_done_pulse) 
                buf_full[rd_sel_reg] <= 1'b0;

            // --- д�����߼� ---
            if (wr_handshake) begin
                if (wr_sel == 0) ram_buf0[wr_ptr] <= s_axis_tdata;
                else             ram_buf1[wr_ptr] <= s_axis_tdata;

                if (wr_finish) begin
                    buf_full[wr_sel] <= 1'b1;         // ��ǵ�ǰ Buffer ��
                    
                    // ��¼����
                    if (wr_sel == 0) len_buf0 <= wr_ptr + 1'b1;
                    else             len_buf1 <= wr_ptr + 1'b1;

                    // �л�
                    wr_sel <= ~wr_sel;
                    wr_ptr <= 0;
                end else begin
                    wr_ptr <= wr_ptr + 1'b1;
                end
            end
        end
    end

    // =========================================================================
    // 3. ��ȡ�߼� (Read Control) - �޸��� Valid ʱ������
    // =========================================================================
    reg [ADDR_WIDTH:0] rd_ptr;
    reg                rd_sel;      // ��ǰ���ڶ��� buffer ����
    reg                rd_active;   // ״̬��־���Ƿ���������ȡ��

    // ��ģ�齻���ź�
    reg  rd_buf_done_pulse; // ֪ͨд����ͷ� Buffer
    reg  rd_sel_reg;        // ��¼�ո��ͷŵ����ĸ� Buffer

    wire [ADDR_WIDTH:0] current_rd_len = (rd_sel == 0) ? len_buf0 : len_buf1;

    // ����߼���ȡ���� (Distributed RAM ģʽ)
    reg [DATA_WIDTH-1:0] ram_rdata_comb;
    always @(*) begin
        if (rd_sel == 0) ram_rdata_comb = ram_buf0[rd_ptr];
        else             ram_rdata_comb = ram_buf1[rd_ptr];
    end

    // ��ȡʹ��������
    // 1. �������� (rd_active) ������ Ready
    // 2. û���У�����ǰ Buffer ���� (buf_full) ��û�����������
    wire rd_enable = (rd_active) ? m_axis_tready : (buf_full[rd_sel] && !rd_buf_done_pulse);

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            rd_ptr            <= 0;
            rd_sel            <= 0;
            rd_active         <= 0;
            rd_buf_done_pulse <= 0;
            rd_sel_reg        <= 0;
            m_axis_tvalid     <= 0;
            m_axis_tdata      <= 0;
            m_axis_tlast      <= 0;
        end else begin
            // �����ź�Ĭ������
            rd_buf_done_pulse <= 0;

            if (rd_enable) begin
                // --- ��һ����ˮ����ַ���� ---
                if (!rd_active) begin
                    // IDLE -> START: ������ȡ
                    rd_active <= 1'b1;
                    rd_ptr    <= 1; // Ԥȡ��һ����ַ
                end else begin
                    // RUNNING: ��ַ����������ж�
                    if (rd_ptr == current_rd_len) begin
                        // ���굱ǰ��
                        rd_active         <= 1'b0;
                        rd_ptr            <= 0;
                        rd_sel            <= ~rd_sel; // �л���ָ��
                        rd_buf_done_pulse <= 1'b1;    // �����ͷ�����
                        rd_sel_reg        <= rd_sel;
                    end else begin
                        rd_ptr <= rd_ptr + 1'b1;
                    end
                end

                // --- �ڶ�����ˮ��������ݴ��� ---
                // ֻҪ���� Active ״̬������������������
                if (rd_active || (buf_full[rd_sel] && !rd_buf_done_pulse)) begin
                    m_axis_tdata  <= ram_rdata_comb;
                    m_axis_tvalid <= 1'b1; // Ĭ�����ߣ�������ݽ�����������

                    // Last �ź��жϣ���ǰָ���� ����-1 (ע��ʱ�����)
                    if (rd_active && (rd_ptr == current_rd_len - 1'b1)) 
                        m_axis_tlast <= 1'b1;
                    else if (!rd_active && (current_rd_len == 1)) 
                        m_axis_tlast <= 1'b1; // �������������Ϊ1
                    else 
                        m_axis_tlast <= 1'b0;

                    // ���޸����ġ������� Last ֮������ Valid
                    // �� rd_ptr ���� current_rd_len ʱ����ʾ��ǰ�������һ�������Ѿ�����һ���ͳ�
                    // ��һ������������״̬�л���
                    if (rd_ptr == current_rd_len) begin
                        // �����һ�� Buffer (buf_full[~rd_sel]) �Ѿ�׼���ã��򱣳� Valid Ϊ 1 (�޷��л�)
                        // �������� Valid�����������Ч����
                        if (buf_full[~rd_sel]) 
                            m_axis_tvalid <= 1'b1; 
                        else 
                            m_axis_tvalid <= 1'b0; 
                    end
                end
            end else if (m_axis_tready) begin
                // ������� Ready ������û������ (rd_enable=0)������ Valid
                m_axis_tvalid <= 1'b0;
                m_axis_tlast  <= 1'b0;
            end
        end
    end

endmodule