`timescale 1ns / 1ps

module tb_shift_ram_buffer;

    // --- 1. �������� ---
    parameter WIDTH = 64;
    parameter DEPTH = 256;

    // --- 2. �źŶ��� ---
    reg clk;
    reg ce;
    reg [WIDTH-1:0] d;
    wire [WIDTH-1:0] q;

    // --- 3. ʵ���� DUT ---
    shift_ram_buffer_counter #(
        .WIDTH(WIDTH),
        .DEPTH(DEPTH)
    ) u_dut (
        .clk(clk),
        .ce(ce),
        .d(d),
        .q(q)
    );

    // --- 4. ʱ������ ---
    initial begin
        clk = 0;
        forever #5 clk = ~clk; // 100MHz
    end

    // --- 5. �����߼� ---
    integer i;
    reg [WIDTH-1:0] expected_value;
    
    initial begin
        // ��ʼ��
        ce = 0;
        d = 0;
        
        #20;
        $display("��ʼ���� shift_ram_buffer");
        $display("WIDTH=%0d, DEPTH=%0d", WIDTH, DEPTH);
        
        // === ���� 1: �����ݲ��� ===
        $display("\n[����1] ������������");
        ce = 1;
        
        for (i = 0; i < 10; i = i + 1) begin
            d = i + 100; // ���ݣ�100, 101, 102...
            @(posedge clk);
            $display("ʱ�� %0t: ����=%h, ���=%h", $time, d, q);
        end
        
        // === ���� 2: ��Ȳ��� ===
        $display("\n[����2] ��������ӳ�");
        
        // ����һ������ֵ��Ȼ��ȴ�DEPTH�����ڿ����
        d = 64'hDEADBEEF;
        @(posedge clk);
        
        ce = 0; // ��ͣ����
        d = 0;
        
        // �ȴ�DEPTH������
        repeat(DEPTH) @(posedge clk);
        
        ce = 1;
        if (q === 64'hDEADBEEF) begin
            $display("��Ȳ���ͨ��: �ӳ�%0d�����ں������ȷ", DEPTH);
        end else begin
            $display("��Ȳ���ʧ��: ����=DEADBEEF, ʵ��=%h", q);
        end
        
        // === ���� 3: ce�źſ��Ʋ��� ===
        $display("\n[����3] ����ce�źſ���");
        
        for (i = 0; i < 20; i = i + 1) begin
            // ÿ��һ������ʹ��һ��
            ce = (i % 2 == 0);
            d = i + 200;
            @(posedge clk);
            if (ce) begin
                $display("ʱ�� %0t: ce=1, ����=%h, ���=%h", $time, d, q);
            end
        end
        
        // === ���� 4: ���Ʋ��� ===
        $display("\n[����4] ����ָ�뻷��");
        ce = 1;
        
        // ���ͳ���DEPTH������
        for (i = 0; i < DEPTH + 10; i = i + 1) begin
            d = i + 300;
            @(posedge clk);
            if (i >= DEPTH) begin
                $display("ʱ�� %0t: ����=%h, ���=%h (�ѻ���)", $time, d, q);
            end
        end
        
        ce = 0;
        #50;
        
        $display("\n�������");
        $finish;
    end

endmodule