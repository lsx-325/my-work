// `timescale 1ns / 1ps

// module fpga_top_level #(
//     parameter AXIS_DATA_WIDTH = 64,      // AXI Stream λ��
//     parameter NUM_IN_CHANNELS = 8,       // ����ͨ�����ж�
//     parameter DATA_WIDTH      = 8,       // ����/Ȩ��λ��
//     parameter ACCUM_WIDTH     = 32,      // �ۼ�λ��
//     parameter FILTER_SIZE     = 3,       // 3x3 ���
//     parameter IMG_WIDTH       = 256,     // ͼ����
//     parameter IMG_HEIGHT      = 256,     // ͼ��߶�
//     parameter BRAM_DEPTH      = 512      // Ȩ�� BRAM ���
// )(
//     input                                   clk,
//     input                                   rst_n,

//     // 1. ͼ������ (AXI-Stream)
//     input                                   s_axis_img_tvalid,
//     output                                  s_axis_img_tready,
//     input      [AXIS_DATA_WIDTH-1:0]        s_axis_img_tdata,
//     input                                   s_axis_img_tlast,

//     // 2. Ȩ������ (AXI-Stream) - �㲥������ BRAM
//     input                                   s_axis_w_tvalid,
//     output reg                              s_axis_w_tready,
//     input      [AXIS_DATA_WIDTH-1:0]        s_axis_w_tdata,
//     input                                   s_axis_w_tlast,

//     // 3. ������ (AXI-Stream)
//     output                                  m_axis_res_tvalid,
//     input                                   m_axis_res_tready,
//     output     [AXIS_DATA_WIDTH-1:0]        m_axis_res_tdata,
//     output     [AXIS_DATA_WIDTH/8-1:0]      m_axis_res_tkeep,
//     output                                  m_axis_res_tlast,

//     // 4. ����������
//     input                                   i_load_weights,     // Ȩ�ؼ���ʹ��
//     input      [3:0]                        i_target_layer,     // Ȩ�ؼ���Ŀ���/��ID (����ƬѡBRAM)
    
//     input                                   i_start_compute,    // ��ʼ����
    
//     // **��̬Ȩ�ص�ַ����**
//     // ���� PS ��ָ����ǰ����ʹ����һ��Ȩ�� (ʵ������ Batch ���������˲����л�)
//     input      [8:0]                        i_l1_weight_base,   // Layer 1 Ȩ�ػ���ַ
//     input      [8:0]                        i_l2_weight_base,   // Layer 2 Ȩ�ػ���ַ
    
//     output                                  o_compute_done
// );

//     // =========================================================================
//     // ��������
//     // =========================================================================
//     // Layer 1 ��Ҫ��� 8 ��ͨ����ÿ�� Core �� 2 ����������Ҫ 4 �� Core
//     localparam L1_NUM_CORES = 4; 
    
//     // ����λ����
//     localparam WIN_BITS = NUM_IN_CHANNELS * FILTER_SIZE * FILTER_SIZE * DATA_WIDTH;
//     localparam W_BITS   = WIN_BITS; // Ȩ��λ���봰��λ��һ��
//     localparam SUM_BITS = ACCUM_WIDTH + $clog2(NUM_IN_CHANNELS); // 35 bit

//     // =========================================================================
//     // �ڲ��ź�
//     // =========================================================================
    
//     // --- Layer 1 ---
//     wire w_win_valid_1;
//     wire [WIN_BITS-1:0] w_win_1;
    
//     // Layer 1 ���к����ź�����
//     wire [W_BITS-1:0]   w_ka_1 [L1_NUM_CORES-1:0];
//     wire [W_BITS-1:0]   w_kb_1 [L1_NUM_CORES-1:0];
//     wire signed [SUM_BITS-1:0] w_sum_a_1 [L1_NUM_CORES-1:0];
//     wire signed [SUM_BITS-1:0] w_sum_b_1 [L1_NUM_CORES-1:0];
//     wire [L1_NUM_CORES-1:0]    w_valid_1;

//     // ����������� (8 channels * 8 bit = 64 bit)
//     reg  [L1_NUM_CORES*2*DATA_WIDTH-1:0] r_layer1_out_packed; 
//     reg  r_layer1_valid;

//     // --- Layer 2 ---
//     wire w_win_valid_2;
//     wire [WIN_BITS-1:0] w_win_2; // Layer 2 ����Ҳ�� 8 ͨ�� (�� L1 ���ƴ��)
    
//     wire [W_BITS-1:0]   w_ka_2, w_kb_2;
//     wire signed [SUM_BITS-1:0] w_sum_a_2, w_sum_b_2;
//     wire w_valid_2;

//     // --- Ȩ������ ---
//     // ���߼������� BRAM ͬʱ�������ݣ�ͨ��дʹ��(��ַ��λ)����
//     // �����Ϊ��ʼ�� Ready������ Valid �� i_target_layer ����
//     always @(*) s_axis_w_tready = 1'b1;

//     // =========================================================================
//     // 1. Layer 1: Line Buffer (Padding & Window Gen)
//     // =========================================================================
//     line_buffer_with_padding #(
//         .NUM_CHANNELS(NUM_IN_CHANNELS),
//         .DATA_WIDTH  (DATA_WIDTH),
//         .IMG_WIDTH   (IMG_WIDTH),
//         .IMG_HEIGHT  (IMG_HEIGHT)
//     ) u_lb_1 (
//         .clk             (clk),
//         .rst_n           (rst_n),
//         .i_valid         (s_axis_img_tvalid && s_axis_img_tready),
//         .i_data_parallel (s_axis_img_tdata),
//         .o_valid         (w_win_valid_1),
//         .o_windows_packed(w_win_1)
//     );
//     assign s_axis_img_tready = 1'b1; 

//     // =========================================================================
//     // 2. Layer 1: ���м������� (4 Cores -> 8 Output Channels)
//     // =========================================================================
//     genvar i;
//     generate
//         for (i = 0; i < L1_NUM_CORES; i = i + 1) begin : gen_l1_cores
            
//             // 2.1 Ȩ�� BRAM ������ (Bank i)
//             // ÿ�� Core ӵ�ж����� BRAM������˵�� BRAM ��һ���߼�����
//             // ��ַ�߼���Core[i] ��ȡ Base + i
//             weight_bram_controller #(
//                 .BRAM_DEPTH(BRAM_DEPTH)
//             ) u_w_bram_1 (
//                 .clk(clk), .rst_n(rst_n),
//                 // д�˿ڣ����� BRAM ����������
//                 .s_axis_tvalid(s_axis_w_tvalid), 
//                 .s_axis_tready(), // ������ Ready����ֹ��������ͻ������ͳһ����
//                 .s_axis_tdata (s_axis_w_tdata),
//                 .s_axis_tlast (s_axis_w_tlast),
                
//                 // д���ƣ����� target_layer == i ʱ�Ÿ�λд��ַ����ʼ����
//                 // ��������ʵ�ַ�ʱ���أ��ȷ� Core0Ȩ�أ��ٷ� Core1Ȩ��...
//                 .i_write_addr_rst(i_load_weights && (i_target_layer == i)),
                
//                 // �����ƣ���̬��ַ + ƫ��
//                 .i_read_addr(i_l1_weight_base), 
//                 .i_read_en  (1'b1),
                
//                 .o_kernels_A_packed(w_ka_1[i]),
//                 .o_kernels_B_packed(w_kb_1[i])
//             );

//             // 2.2 �������
//             conv_3x3_parallel_top u_conv_1 (
//                 .clk(clk), .rst_n(rst_n),
//                 .i_valid(w_win_valid_1 && i_start_compute),
//                 .i_windows_packed(w_win_1), // ���� Core ������ͬ�����봰��
//                 .i_kernels_A_packed(w_ka_1[i]),
//                 .i_kernels_B_packed(w_kb_1[i]),
//                 .o_final_sum_A(w_sum_a_1[i]),
//                 .o_final_sum_B(w_sum_b_1[i]),
//                 .o_final_valid(w_valid_1[i])
//             );
//         end
//     endgenerate

//     // =========================================================================
//     // 3. Layer 1 -> Layer 2 ������ (ReLU + Quantization + Concatenation)
//     // =========================================================================
//     // ��������
//     function [7:0] quantize;
//         input signed [34:0] val;
//         begin
//             if (val < 0) quantize = 0; // ReLU
//             else if ((val >>> 10) > 255) quantize = 255; // Clip
//             else quantize = val[17:10]; // Scale
//         end
//     endfunction

//     integer j;
//     always @(posedge clk or negedge rst_n) begin
//         if(!rst_n) begin
//             r_layer1_out_packed <= 0;
//             r_layer1_valid <= 0;
//         end else begin
//             // ʹ�� Core 0 �� valid ��Ϊͬ���ź� (�������� Core ͬ��)
//             r_layer1_valid <= w_valid_1[0];
            
//             if (w_valid_1[0]) begin
//                 // ƴ�� 4 �� Core ����� (4 * 2 = 8 Channels)
//                 // Core 0 (Ch 0,1), Core 1 (Ch 2,3), Core 2 (Ch 4,5), Core 3 (Ch 6,7)
//                 // ���� Little-Endian: {Core3_B, Core3_A ... Core0_B, Core0_A}
//                 for (j = 0; j < L1_NUM_CORES; j = j + 1) begin
//                     r_layer1_out_packed[(j*16) +: 8]      <= quantize(w_sum_a_1[j]); // Ch A
//                     r_layer1_out_packed[(j*16 + 8) +: 8]  <= quantize(w_sum_b_1[j]); // Ch B
//                 end
//             end
//         end
//     end

//     // =========================================================================
//     // 4. Layer 2: Line Buffer
//     // =========================================================================
//     // ��ʱ Layer 2 ���յ�����ʵ�� 8 ͨ����������
//     line_buffer_with_padding #(
//         .NUM_CHANNELS(NUM_IN_CHANNELS), // 8
//         .IMG_WIDTH   (IMG_WIDTH),
//         .IMG_HEIGHT  (IMG_HEIGHT)
//     ) u_lb_2 (
//         .clk(clk), .rst_n(rst_n),
//         .i_valid(r_layer1_valid),
//         .i_data_parallel(r_layer1_out_packed),
//         .o_valid(w_win_valid_2),
//         .o_windows_packed(w_win_2)
//     );

//     // =========================================================================
//     // 5. Layer 2: ������� (������ʾ��)
//     // =========================================================================
//     // ���� Layer 2 ֻ��Ҫ��� 2 ��ͨ���� Saver
//     // ��� Layer 2 Ҳ��Ҫ����ͨ��������ͬ��ʹ�� generate ����
    
//     weight_bram_controller #(
//         .BRAM_DEPTH(BRAM_DEPTH)
//     ) u_w_bram_2 (
//         .clk(clk), .rst_n(rst_n),
//         .s_axis_tvalid(s_axis_w_tvalid), 
//         .s_axis_tready(), 
//         .s_axis_tdata (s_axis_w_tdata),
//         .s_axis_tlast (s_axis_w_tlast),
//         // Target ID ��Ϊ 4 (0-3 �� Layer 1 ռ��)
//         .i_write_addr_rst(i_load_weights && (i_target_layer == 4)), 
        
//         .i_read_addr(i_l2_weight_base), // ��̬����ַ
//         .i_read_en  (1'b1),
//         .o_kernels_A_packed(w_ka_2),
//         .o_kernels_B_packed(w_kb_2)
//     );

//     conv_3x3_parallel_top u_conv_2 (
//         .clk(clk), .rst_n(rst_n),
//         .i_valid(w_win_valid_2),
//         .i_windows_packed(w_win_2),
//         .i_kernels_A_packed(w_ka_2),
//         .i_kernels_B_packed(w_kb_2),
//         .o_final_sum_A(w_sum_a_2),
//         .o_final_sum_B(w_sum_b_2),
//         .o_final_valid(w_valid_2)
//     );

//     // =========================================================================
//     // 6. ������
//     // =========================================================================
//     feature_map_saver_axis #(
//         .AXIS_DATA_WIDTH(AXIS_DATA_WIDTH),
//         .INPUT_WIDTH    (ACCUM_WIDTH + $clog2(NUM_IN_CHANNELS)), 
//         .OUTPUT_WIDTH   (8),
//         .QUANT_SHIFT    (10)
//     ) u_saver (
//         .clk           (clk),
//         .rst_n         (rst_n),
//         .i_valid       (w_valid_2),
//         .i_data_A      (w_sum_a_2),
//         .i_data_B      (w_sum_b_2),
//         .i_total_pixels(IMG_WIDTH * IMG_HEIGHT),
        
//         .m_axis_tvalid (m_axis_res_tvalid),
//         .m_axis_tready (m_axis_res_tready),
//         .m_axis_tdata  (m_axis_res_tdata),
//         .m_axis_tkeep  (m_axis_res_tkeep),
//         .m_axis_tlast  (m_axis_res_tlast)
//     );
    
//     assign o_compute_done = m_axis_res_tvalid && m_axis_res_tlast;

// endmodule
`timescale 1ns / 1ps

module fpga_top_level #(
    parameter AXIS_DATA_WIDTH = 64,      // AXI Stream λ�� (8ͨ�� * 8bit)
    parameter NUM_IN_CHANNELS = 8,       // ����ͨ�����ж�
    parameter DATA_WIDTH      = 8,       // ����/Ȩ��λ��
    parameter ACCUM_WIDTH     = 32,      // �ۼ�λ��
    parameter FILTER_SIZE     = 3,       // 3x3 ���
    parameter IMG_WIDTH       = 256,     // ͼ����
    parameter IMG_HEIGHT      = 256,     // ͼ��߶�
    parameter BRAM_DEPTH      = 512      // Ȩ�� BRAM ���
)(
    input                                   clk,
    input                                   rst_n,

    // 1. ͼ������ (AXI-Stream)
    input                                   s_axis_img_tvalid,
    output                                  s_axis_img_tready, // ���޸ġ������� PingPong ����
    input      [AXIS_DATA_WIDTH-1:0]        s_axis_img_tdata,
    input                                   s_axis_img_tlast,

    // 2. Ȩ������ (AXI-Stream) - �㲥������ BRAM
    input                                   s_axis_w_tvalid,
    output                                  s_axis_w_tready,
    input      [AXIS_DATA_WIDTH-1:0]        s_axis_w_tdata,
    input                                   s_axis_w_tlast,

    // 3. ������ (AXI-Stream)
    output                                  m_axis_res_tvalid,
    input                                   m_axis_res_tready,
    output     [AXIS_DATA_WIDTH-1:0]        m_axis_res_tdata,
    output     [AXIS_DATA_WIDTH/8-1:0]      m_axis_res_tkeep,
    output                                  m_axis_res_tlast,

    // 4. ����������
    input                                   i_load_weights,     // Ȩ�ؼ���ʹ��
    input      [3:0]                        i_target_layer,     // Ȩ�ؼ���Ŀ���ID
    input                                   i_start_compute,    // ��ʼ����
    
    // **��̬Ȩ�ص�ַ����**
    input      [8:0]                        i_l1_weight_base,   
    input      [8:0]                        i_l2_weight_base, 
    
    output                                  o_compute_done
);

    // =========================================================================
    // ��������
    // =========================================================================
    localparam L1_NUM_CORES = 4;
    // ����λ����
    localparam WIN_BITS = NUM_IN_CHANNELS * FILTER_SIZE * FILTER_SIZE * DATA_WIDTH;
    localparam W_BITS   = WIN_BITS; 
    localparam SUM_BITS = ACCUM_WIDTH + $clog2(NUM_IN_CHANNELS);

    // =========================================================================
    // �ڲ��ź�
    // =========================================================================
    
    // --- Layer 1 ---
    wire w_win_valid_1;
    wire [WIN_BITS-1:0] w_win_1;
    
    wire [W_BITS-1:0]   w_ka_1 [L1_NUM_CORES-1:0];
    wire [W_BITS-1:0]   w_kb_1 [L1_NUM_CORES-1:0];
    wire signed [SUM_BITS-1:0] w_sum_a_1 [L1_NUM_CORES-1:0];
    wire signed [SUM_BITS-1:0] w_sum_b_1 [L1_NUM_CORES-1:0];
    wire [L1_NUM_CORES-1:0]    w_valid_1;

    // �����������
    reg  [L1_NUM_CORES*2*DATA_WIDTH-1:0] r_layer1_out_packed;
    reg  r_layer1_valid;

    // --- Layer 2 ---
    wire w_win_valid_2;
    wire [WIN_BITS-1:0] w_win_2;
    wire w_l2_ready; // Layer 2 �� PingPong ��ѹ�ź� (�����ݲ����� L1 ��ͣ)
    
    wire [W_BITS-1:0]   w_ka_2, w_kb_2;
    wire signed [SUM_BITS-1:0] w_sum_a_2, w_sum_b_2;
    wire w_valid_2;

    // Ȩ�� Ready �ź�Ĭ������
    assign s_axis_w_tready = 1'b1;

    // =========================================================================
    // 1. Layer 1: ���뻺��ϵͳ (PingPong + Padding + Window Gen)
    // =========================================================================
    // ���޸ġ��滻ԭ�е� line_buffer_with_padding
    
    system_top u_sys_top_l1 (
        .sys_clk        (clk),
        .sys_rst_n      (rst_n),
        
        // �ⲿ DMA / AXIS ����
        .dma_valid      (s_axis_img_tvalid),
        .dma_data       (s_axis_img_tdata),
        .dma_ready      (s_axis_img_tready), // �����ѹ�źŸ��ⲿ AXI
        
        // ��̬���� (ʹ�� Parameter ת��)
        .cfg_width      (IMG_WIDTH[15:0]),
        .cfg_height     (IMG_HEIGHT[15:0]),
        .cfg_pad_en     (1'b1), // Layer 1 ���� Padding (Same)
        
        // ����� Layer 1 �����
        .conv_valid     (w_win_valid_1),
        .conv_window    (w_win_1)
    );

    // =========================================================================
    // 2. Layer 1: ���м������� (4 Cores -> 8 Output Channels)
    // =========================================================================
    genvar i;
    generate
        for (i = 0; i < L1_NUM_CORES; i = i + 1) begin : gen_l1_cores
            
            // 2.1 Ȩ�� BRAM
            weight_bram_controller #(.BRAM_DEPTH(BRAM_DEPTH)) u_w_bram_1 (
                .clk(clk), .rst_n(rst_n),
                .s_axis_tvalid(s_axis_w_tvalid), 
                .s_axis_tready(), 
                .s_axis_tdata (s_axis_w_tdata),
                .s_axis_tlast (s_axis_w_tlast),
                .i_write_addr_rst(i_load_weights && (i_target_layer == i)),
                .i_read_addr(i_l1_weight_base), 
                .i_read_en  (1'b1),
                .o_kernels_A_packed(w_ka_1[i]),
                .o_kernels_B_packed(w_kb_1[i])
            );

            // 2.2 �������
            // ע�⣺start_compute ������Ч��
            conv_3x3_parallel_top u_conv_1 (
                .clk(clk), .rst_n(rst_n),
                .i_valid(w_win_valid_1 && i_start_compute),
                .i_windows_packed(w_win_1), 
                .i_kernels_A_packed(w_ka_1[i]),
                .i_kernels_B_packed(w_kb_1[i]),
                .o_final_sum_A(w_sum_a_1[i]),
                .o_final_sum_B(w_sum_b_1[i]),
                .o_final_valid(w_valid_1[i])
            );
        end
    endgenerate

    // =========================================================================
    // 3. Layer 1 -> Layer 2 ������ (ReLU + Quantization)
    // =========================================================================
    function [7:0] quantize;
        input signed [34:0] val;
        begin
            if (val < 0) quantize = 0;                   // ReLU
            else if ((val >>> 10) > 255) quantize = 255; // Clip
            else quantize = val[17:10];                  // Scale
        end
    endfunction

    integer j;
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            r_layer1_out_packed <= 0;
            r_layer1_valid <= 0;
        end else begin
            // ���߼����������� Core ͬ�����
            r_layer1_valid <= w_valid_1[0];
            
            if (w_valid_1[0]) begin
                for (j = 0; j < L1_NUM_CORES; j = j + 1) begin
                    r_layer1_out_packed[(j*16) +: 8]      <= quantize(w_sum_a_1[j]);
                    r_layer1_out_packed[(j*16 + 8) +: 8]  <= quantize(w_sum_b_1[j]);
                end
            end
        end
    end

    // =========================================================================
    // 4. Layer 2: ���뻺��ϵͳ (PingPong + Padding)
    // =========================================================================
    // ���޸ġ��滻ԭ�е� line_buffer_with_padding
    // Layer 1 �������� (8ͨ��, 64bit) ���� Layer 2 �� Ping-Pong Buffer
    
    system_top u_sys_top_l2 (
        .sys_clk        (clk),
        .sys_rst_n      (rst_n),
        
        // �������� Layer 1 ������
        .dma_valid      (r_layer1_valid),
        .dma_data       (r_layer1_out_packed),
        .dma_ready      (w_l2_ready), // ����� Ready ������������أ����������Ҫ�����ӵĿ���
                                      // ���������Ӧ������ Layer 1 ��ͣ��ˮ��
                                      
        // ��̬���� (Layer 2 �ߴ��� Layer 1 ��ͬ)
        .cfg_width      (IMG_WIDTH[15:0]),
        .cfg_height     (IMG_HEIGHT[15:0]),
        .cfg_pad_en     (1'b1), // Layer 2 ͬ������ Padding
        
        // ����� Layer 2 �����
        .conv_valid     (w_win_valid_2),
        .conv_window    (w_win_2)
    );

    // =========================================================================
    // 5. Layer 2: �������
    // =========================================================================
    weight_bram_controller #(.BRAM_DEPTH(BRAM_DEPTH)) u_w_bram_2 (
        .clk(clk), .rst_n(rst_n),
        .s_axis_tvalid(s_axis_w_tvalid), 
        .s_axis_tready(), 
        .s_axis_tdata (s_axis_w_tdata),
        .s_axis_tlast (s_axis_w_tlast),
        .i_write_addr_rst(i_load_weights && (i_target_layer == 4)), 
        .i_read_addr(i_l2_weight_base), 
        .i_read_en  (1'b1),
        .o_kernels_A_packed(w_ka_2),
        .o_kernels_B_packed(w_kb_2)
    );

    conv_3x3_parallel_top u_conv_2 (
        .clk(clk), .rst_n(rst_n),
        .i_valid(w_win_valid_2),
        .i_windows_packed(w_win_2),
        .i_kernels_A_packed(w_ka_2),
        .i_kernels_B_packed(w_kb_2),
        .o_final_sum_A(w_sum_a_2),
        .o_final_sum_B(w_sum_b_2),
        .o_final_valid(w_valid_2)
    );

    // =========================================================================
    // 6. ������
    // =========================================================================
    feature_map_saver_axis #(
        .AXIS_DATA_WIDTH(AXIS_DATA_WIDTH),
        .INPUT_WIDTH    (ACCUM_WIDTH + $clog2(NUM_IN_CHANNELS)), 
        .OUTPUT_WIDTH   (8),
        .QUANT_SHIFT    (10)
    ) u_saver (
        .clk           (clk),
        .rst_n         (rst_n),
        .i_valid       (w_valid_2),
        .i_data_A      (w_sum_a_2),
        .i_data_B      (w_sum_b_2),
        .i_total_pixels(IMG_WIDTH * IMG_HEIGHT),
        .m_axis_tvalid (m_axis_res_tvalid),
        .m_axis_tready (m_axis_res_tready),
        .m_axis_tdata  (m_axis_res_tdata),
        .m_axis_tkeep  (m_axis_res_tkeep),
        .m_axis_tlast  (m_axis_res_tlast)
    );

    assign o_compute_done = m_axis_res_tvalid && m_axis_res_tlast;

endmodule