//module dsp2x8 (                                         // ����8bit�˷�����һ��DSP,���λ��15λ
//    input                   clk  ,
//    input                   rst_n,
//    input                   CE   ,
//    input  signed [8-1:0]   D    ,
//    input  signed [8-1:0]   WA   ,
//    input  signed [8-1:0]   WB   ,
//    output        [15-1:0]    QA   ,
//    output        [15-1:0]    QB
//);
    
//    reg  signed [23:0] w;
//    reg  signed [7:0]  d_r;
//    (* use_dsp="yes" *)
//    reg  signed [32:0] res;
//    wire signed [16-1:0] qb;
//    reg  ce_r;
    
//    assign QA = (^res[15:14])? 15'd16383: res[14:0];
//    assign QB = (^qb[15:14])? 15'd16383: qb[14:0];
//    assign qb = res[31:16] + res[15]; 

//    always @ (posedge clk)
//        if (!rst_n)
//            ce_r <= 'b0;
//        else
//            ce_r <= CE;
    
//    always @ (posedge clk)
//        if (CE) begin
//            d_r <= D;
//            w   <= WA + (WB <<< 16);
//        end
        
//    always @ (posedge clk)
//        if (ce_r)
//            res <= d_r * w;
            
//endmodule
//// ����ģ��
///*
//    dsp2x8 dsp2x8_u (
//        .clk  (clk  ), // input
//        .CE   (CE   ), // input                
//        .D    (D    ), // input  signed [7:0]  
//        .WA   (WA   ), // input  signed [7:0]  
//        .WB   (WB   ), // input  signed [7:0]
//        .QA   (QA   ), // output        [15:0] 
//        .QB   (QB   )  // output        [15:0] 
//    );
//*/
module dsp2x8 (                        //// ����8bit�˷�����һ��DSP,���λ��16λ                         
    input                  clk  ,
    input                  rst_n,
    input                  CE   ,
    input  signed [7:0]    D    ,
    input  signed [7:0]    WA   ,
    input  signed [7:0]    WB   ,
    output signed [15:0]   QA   , // �޸ĵ�1�����λ���Ϊ 16 bit
    output signed [15:0]   QB     // �޸ĵ�1�����λ���Ϊ 16 bit
);

    // �޸ĵ�2�������޸���w ��չΪ 25 bit
    // 25 bit ��Χ��-16,777,216 �� +16,777,215
    // �������� (-128 << 16) + (-1) = -8,388,609���������Ϊ����
    reg  signed [24:0] w;     
    
    reg  signed [7:0]  d_r;
    
    // 33 bit (8 bit * 25 bit) �պ����� DSP48
    (* use_dsp="yes" *)
    reg  signed [32:0] res;   
    
    wire signed [15:0] qb_wire; // �ڲ� wire Ҳ��Ϊ 16 bit
    reg  ce_r;

    // �޸ĵ�3���Ƴ� 15-bit ���ͽض��߼�
    // ��� QA/QB �� 16-bit�������ֱ������������� res[15:14] �����
    assign QA = res[15:0]; 
    assign QB = qb_wire;

    // ��λ��ȡ�߼����ֲ��䣺
    // ʹ�� res[15] (��λ���ֵķ���λ) ��������λ
    assign qb_wire = res[31:16] + res[15];

    always @ (posedge clk)
        if (!rst_n)
            ce_r <= 'b0;
        else
            ce_r <= CE;

    always @ (posedge clk)
        if (CE) begin
            d_r <= D;
            // �޸ĵ�2ԭ��
            // WB(8bit) ���� 16 λ��Verilog ���Զ������� 25-bit ������������
            // �ܹ���ȷ�������λ��λ
            w   <= WA + (WB <<< 16);
        end
        
    always @ (posedge clk)
        if (ce_r)
            res <= d_r * w; 

endmodule